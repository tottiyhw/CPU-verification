module CU_module(clr,clk,Op,IRFunc,IRFunc1,IRFunc2,zero,OV,lt,gt,LLbit,fp,IR,TrapAddr,CtrlA,CtrlALUOut,CtrlB,CtrlCP0,CtrlCP0_ASID,CtrlCP0_EPC,CtrlCP0_ExCode,CtrlCP1,CtrlConditionReg,CtrlDMem,CtrlDR,CtrlDR0,CtrlGPR,CtrlHi,CtrlIR,CtrlLLbit,CtrlLo,CtrlOVReg,CtrlPC,CtrlPCInc,CtrlPIDReg,CtrlMux1_1,CtrlMux1_2,CtrlMux1_3,CtrlMux1_4,CtrlMux1_5,CtrlMux2_1,CtrlMux3_1,CtrlMux4_1,CtrlMux5_1,CtrlMux6_1,CtrlMux7_1,CtrlMux7_2,CtrlMux9_1,CtrlMux10_1,CtrlMux10_2,CtrlMux11_1,CtrlMux12_1,CtrlMux12_2,CtrlMux12_3,CtrlMux12_4,CtrlMux12_5,CtrlMux12_6,CtrlMux12_7,CtrlMux12_8,CtrlMux12_9,CtrlMux12_10,CtrlMux12_11,CtrlMux13_1,CtrlMux13_2,CtrlMux13_3,CtrlMux14_1,CtrlMux14_2,CtrlMux15_1,CtrlMux15_2,CtrlMux15_3,CtrlMux16_1,CtrlMux16_2,CtrlMux16_3,CtrlMux17_1,CtrlMux17_2,CtrlMux18_1,CtrlMux18_2,CtrlMux18_3,CtrlMux18_4,CtrlMux18_5,CtrlMux18_6,CtrlMux18_7,CtrlMux18_8,CtrlMux18_9,CtrlMux19_1,CtrlMux19_2,CtrlMux20_1,CtrlMux21_1,CtrlMux22_1,CtrlMux23_1,CtrlMux24_1,CtrlMux25_1,CtrlMux26_1,CtrlMux26_2,CtrlMux27_1,CtrlMux28_1,CtrlMux28_2,CtrlMux29_1,CtrlMux29_2,CtrlMux30_1,CtrlMux31_1,CtrlMux31_2,CtrlMux31_3,CtrlMux32_1,CtrlMux33_1,CtrlMux33_2,CtrlMux34_1,CtrlMux34_2,CtrlMux35_1,CtrlMux36_1,CtrlMux37_1,CtrlMux38_1,CtrlMux38_2,CtrlMux38_3,CtrlMux38_4,CtrlMux38_5,CtrlMux38_6,CtrlMux38_7,CtrlMux38_8,CtrlMux39_1,CtrlMux40_1,CtrlMux41_1,CtrlMux41_2,CtrlMux41_3,CtrlMux41_4,CtrlMux41_5,CtrlMux41_6,CtrlMux41_7,CtrlMux41_8,CtrlMux41_9,CtrlMux41_10,CtrlMux41_11,CtrlMux42_1,CtrlMux43_1,CtrlMux44_1,CtrlMux44_2,CtrlMux45_1,CtrlMux46_1,CtrlMux46_2,CtrlMux46_3,CtrlMux46_4,CtrlMux47_1,CtrlMux48_1,CtrlMux49_1,CtrlMux49_2,CtrlMux49_3,CtrlMux50_1,CtrlMux50_2,CtrlMux51_1,CtrlMux51_2,CtrlMux52_1,CtrlMux53_1,CtrlMux53_2,CtrlMux54_1,CtrlMux55_1,CtrlMux56_1,CtrlMux57_1,CtrlMux58_1,CtrlMux59_1,CtrlMux60_1,CtrlMux61_1,CtrlMux64_1,CtrlMux65_1,CtrlMux68_1,CtrlMux69_1,CtrlMux70_1,CtrlMux71_1,CtrlMux72_1);
input clr;
input clk;
input [5:0]Op;
input [5:0]IRFunc;
input [4:0]IRFunc1;
input [4:0]IRFunc2;
input zero;
input OV;
input lt;
input gt;
input LLbit;
input fp;
input [31:0]IR;
output [31:0]TrapAddr;
output CtrlA;
output CtrlALUOut;
output CtrlB;
output CtrlCP0;
output CtrlCP0_ASID;
output CtrlCP0_EPC;
output CtrlCP0_ExCode;
output CtrlCP1;
output CtrlConditionReg;
output CtrlDMem;
output CtrlDR;
output CtrlDR0;
output CtrlGPR;
output CtrlHi;
output CtrlIR;
output CtrlLLbit;
output CtrlLo;
output CtrlOVReg;
output CtrlPC;
output CtrlPCInc;
output CtrlPIDReg;
output CtrlMux1_1;
output CtrlMux1_2;
output CtrlMux1_3;
output CtrlMux1_4;
output CtrlMux1_5;
output CtrlMux2_1;
output CtrlMux3_1;
output CtrlMux4_1;
output CtrlMux5_1;
output CtrlMux6_1;
output CtrlMux7_1;
output CtrlMux7_2;
output CtrlMux9_1;
output CtrlMux10_1;
output CtrlMux10_2;
output CtrlMux11_1;
output CtrlMux12_1;
output CtrlMux12_2;
output CtrlMux12_3;
output CtrlMux12_4;
output CtrlMux12_5;
output CtrlMux12_6;
output CtrlMux12_7;
output CtrlMux12_8;
output CtrlMux12_9;
output CtrlMux12_10;
output CtrlMux12_11;
output CtrlMux13_1;
output CtrlMux13_2;
output CtrlMux13_3;
output CtrlMux14_1;
output CtrlMux14_2;
output CtrlMux15_1;
output CtrlMux15_2;
output CtrlMux15_3;
output CtrlMux16_1;
output CtrlMux16_2;
output CtrlMux16_3;
output CtrlMux17_1;
output CtrlMux17_2;
output CtrlMux18_1;
output CtrlMux18_2;
output CtrlMux18_3;
output CtrlMux18_4;
output CtrlMux18_5;
output CtrlMux18_6;
output CtrlMux18_7;
output CtrlMux18_8;
output CtrlMux18_9;
output CtrlMux19_1;
output CtrlMux19_2;
output CtrlMux20_1;
output CtrlMux21_1;
output CtrlMux22_1;
output CtrlMux23_1;
output CtrlMux24_1;
output CtrlMux25_1;
output CtrlMux26_1;
output CtrlMux26_2;
output CtrlMux27_1;
output CtrlMux28_1;
output CtrlMux28_2;
output CtrlMux29_1;
output CtrlMux29_2;
output CtrlMux30_1;
output CtrlMux31_1;
output CtrlMux31_2;
output CtrlMux31_3;
output CtrlMux32_1;
output CtrlMux33_1;
output CtrlMux33_2;
output CtrlMux34_1;
output CtrlMux34_2;
output CtrlMux35_1;
output CtrlMux36_1;
output CtrlMux37_1;
output CtrlMux38_1;
output CtrlMux38_2;
output CtrlMux38_3;
output CtrlMux38_4;
output CtrlMux38_5;
output CtrlMux38_6;
output CtrlMux38_7;
output CtrlMux38_8;
output CtrlMux39_1;
output CtrlMux40_1;
output CtrlMux41_1;
output CtrlMux41_2;
output CtrlMux41_3;
output CtrlMux41_4;
output CtrlMux41_5;
output CtrlMux41_6;
output CtrlMux41_7;
output CtrlMux41_8;
output CtrlMux41_9;
output CtrlMux41_10;
output CtrlMux41_11;
output CtrlMux42_1;
output CtrlMux43_1;
output CtrlMux44_1;
output CtrlMux44_2;
output CtrlMux45_1;
output CtrlMux46_1;
output CtrlMux46_2;
output CtrlMux46_3;
output CtrlMux46_4;
output CtrlMux47_1;
output CtrlMux48_1;
output CtrlMux49_1;
output CtrlMux49_2;
output CtrlMux49_3;
output CtrlMux50_1;
output CtrlMux50_2;
output CtrlMux51_1;
output CtrlMux51_2;
output CtrlMux52_1;
output CtrlMux53_1;
output CtrlMux53_2;
output CtrlMux54_1;
output CtrlMux55_1;
output CtrlMux56_1;
output CtrlMux57_1;
output CtrlMux58_1;
output CtrlMux59_1;
output CtrlMux60_1;
output CtrlMux61_1;
output CtrlMux64_1;
output CtrlMux65_1;
output CtrlMux68_1;
output CtrlMux69_1;
output CtrlMux70_1;
output CtrlMux71_1;
output CtrlMux72_1;
wire P0,P1,P2,P3,P4,Reset;
wire CtrlFunc00;
wire CtrlFunc01;
wire CtrlFunc02;
wire CtrlFunc03;
wire CtrlFunc04;
wire CtrlFunc05;
wire CtrlFunc06;
wire CtrlFunc07;
wire CtrlFunc08;
wire CtrlFunc09;
wire CtrlFunc0a;
wire CtrlFunc0b;
wire CtrlFunc0c;
wire CtrlFunc0d;
wire CtrlFunc10;
wire CtrlFunc101;
wire CtrlFunc108;
wire CtrlFunc109;
wire CtrlFunc10a;
wire CtrlFunc10b;
wire CtrlFunc10c;
wire CtrlFunc10e;
wire CtrlFunc11;
wire CtrlFunc110;
wire CtrlFunc111;
wire CtrlFunc12;
wire CtrlFunc13;
wire CtrlFunc18;
wire CtrlFunc19;
wire CtrlFunc1a;
wire CtrlFunc1b;
wire CtrlFunc20;
wire CtrlFunc200;
wire CtrlFunc204;
wire CtrlFunc208;
wire CtrlFunc21;
wire CtrlFunc22;
wire CtrlFunc23;
wire CtrlFunc24;
wire CtrlFunc25;
wire CtrlFunc26;
wire CtrlFunc27;
wire CtrlFunc2a;
wire CtrlFunc2b;
wire CtrlFunc30;
wire CtrlFunc31;
wire CtrlFunc32;
wire CtrlFunc33;
wire CtrlFunc34;
wire CtrlFunc36;
wire CtrlOP00;
wire CtrlOP01;
wire CtrlOP02;
wire CtrlOP03;
wire CtrlOP04;
wire CtrlOP05;
wire CtrlOP06;
wire CtrlOP07;
wire CtrlOP08;
wire CtrlOP09;
wire CtrlOP0a;
wire CtrlOP0b;
wire CtrlOP0c;
wire CtrlOP0d;
wire CtrlOP0e;
wire CtrlOP0f;
wire CtrlOP10;
wire CtrlOP11;
wire CtrlOP1c;
wire CtrlOP20;
wire CtrlOP21;
wire CtrlOP22;
wire CtrlOP23;
wire CtrlOP24;
wire CtrlOP25;
wire CtrlOP26;
wire CtrlOP28;
wire CtrlOP29;
wire CtrlOP2a;
wire CtrlOP2b;
wire CtrlOP2e;
wire CtrlOP30;
wire CtrlOP38;
Initial_model Initial(.clr(clr),.clk(clk),.P0(P0),.P1(P1),.P2(P2),.P3(P3),.P4(P4),.Reset(Reset),.Op(Op),.IRFunc(IRFunc),.IRFunc1(IRFunc1),.IRFunc2(IRFunc2),.IR(IR),.nop(nop),.TrapAddr(TrapAddr),.CtrlFunc00(CtrlFunc00),.CtrlFunc01(CtrlFunc01),.CtrlFunc02(CtrlFunc02),.CtrlFunc03(CtrlFunc03),.CtrlFunc04(CtrlFunc04),.CtrlFunc05(CtrlFunc05),.CtrlFunc06(CtrlFunc06),.CtrlFunc07(CtrlFunc07),.CtrlFunc08(CtrlFunc08),.CtrlFunc09(CtrlFunc09),.CtrlFunc0a(CtrlFunc0a),.CtrlFunc0b(CtrlFunc0b),.CtrlFunc0c(CtrlFunc0c),.CtrlFunc0d(CtrlFunc0d),.CtrlFunc10(CtrlFunc10),.CtrlFunc101(CtrlFunc101),.CtrlFunc108(CtrlFunc108),.CtrlFunc109(CtrlFunc109),.CtrlFunc10a(CtrlFunc10a),.CtrlFunc10b(CtrlFunc10b),.CtrlFunc10c(CtrlFunc10c),.CtrlFunc10e(CtrlFunc10e),.CtrlFunc11(CtrlFunc11),.CtrlFunc110(CtrlFunc110),.CtrlFunc111(CtrlFunc111),.CtrlFunc12(CtrlFunc12),.CtrlFunc13(CtrlFunc13),.CtrlFunc18(CtrlFunc18),.CtrlFunc19(CtrlFunc19),.CtrlFunc1a(CtrlFunc1a),.CtrlFunc1b(CtrlFunc1b),.CtrlFunc20(CtrlFunc20),.CtrlFunc200(CtrlFunc200),.CtrlFunc204(CtrlFunc204),.CtrlFunc208(CtrlFunc208),.CtrlFunc21(CtrlFunc21),.CtrlFunc22(CtrlFunc22),.CtrlFunc23(CtrlFunc23),.CtrlFunc24(CtrlFunc24),.CtrlFunc25(CtrlFunc25),.CtrlFunc26(CtrlFunc26),.CtrlFunc27(CtrlFunc27),.CtrlFunc2a(CtrlFunc2a),.CtrlFunc2b(CtrlFunc2b),.CtrlFunc30(CtrlFunc30),.CtrlFunc31(CtrlFunc31),.CtrlFunc32(CtrlFunc32),.CtrlFunc33(CtrlFunc33),.CtrlFunc34(CtrlFunc34),.CtrlFunc36(CtrlFunc36),.CtrlOP00(CtrlOP00),.CtrlOP01(CtrlOP01),.CtrlOP02(CtrlOP02),.CtrlOP03(CtrlOP03),.CtrlOP04(CtrlOP04),.CtrlOP05(CtrlOP05),.CtrlOP06(CtrlOP06),.CtrlOP07(CtrlOP07),.CtrlOP08(CtrlOP08),.CtrlOP09(CtrlOP09),.CtrlOP0a(CtrlOP0a),.CtrlOP0b(CtrlOP0b),.CtrlOP0c(CtrlOP0c),.CtrlOP0d(CtrlOP0d),.CtrlOP0e(CtrlOP0e),.CtrlOP0f(CtrlOP0f),.CtrlOP10(CtrlOP10),.CtrlOP11(CtrlOP11),.CtrlOP1c(CtrlOP1c),.CtrlOP20(CtrlOP20),.CtrlOP21(CtrlOP21),.CtrlOP22(CtrlOP22),.CtrlOP23(CtrlOP23),.CtrlOP24(CtrlOP24),.CtrlOP25(CtrlOP25),.CtrlOP26(CtrlOP26),.CtrlOP28(CtrlOP28),.CtrlOP29(CtrlOP29),.CtrlOP2a(CtrlOP2a),.CtrlOP2b(CtrlOP2b),.CtrlOP2e(CtrlOP2e),.CtrlOP30(CtrlOP30),.CtrlOP38(CtrlOP38));
assign CtrlA=(P1&CtrlOP00&CtrlFunc20)|(P1&CtrlOP00&CtrlFunc22)|(P1&CtrlOP00&CtrlFunc21)|(P1&CtrlOP00&CtrlFunc23)|(P1&CtrlOP00&CtrlFunc24)|(P1&CtrlOP00&CtrlFunc25)|(P1&CtrlOP00&CtrlFunc26)|(P1&CtrlOP00&CtrlFunc27)|(P1&CtrlOP00&CtrlFunc2a)|(P1&CtrlOP00&CtrlFunc2b)|(P1&CtrlOP08)|(P1&CtrlOP09)|(P1&CtrlOP0a)|(P1&CtrlOP0b)|(P1&CtrlOP0c)|(P1&CtrlOP0d)|(P1&CtrlOP0e)|(P1&CtrlOP00&CtrlFunc04)|(P1&CtrlOP00&CtrlFunc06)|(P1&CtrlOP00&CtrlFunc07)|(P1&CtrlOP00&CtrlFunc18)|(P1&CtrlOP00&CtrlFunc19)|(P1&CtrlOP00&CtrlFunc1a)|(P1&CtrlOP00&CtrlFunc1b)|(P1&CtrlOP1c&CtrlFunc02)|(P1&CtrlOP04)|(P1&CtrlOP05)|(P1&CtrlOP07)|(P1&CtrlOP06)|(P1&CtrlOP01)|(P1&CtrlOP01&CtrlFunc101)|(P1&CtrlOP01&CtrlFunc110)|(P1&CtrlOP01&CtrlFunc111)|(P1&CtrlOP00&CtrlFunc30)|(P1&CtrlOP00&CtrlFunc31)|(P1&CtrlOP00&CtrlFunc32)|(P1&CtrlOP00&CtrlFunc33)|(P1&CtrlOP00&CtrlFunc34)|(P1&CtrlOP00&CtrlFunc36)|(P1&CtrlOP01&CtrlFunc108)|(P1&CtrlOP01&CtrlFunc109)|(P1&CtrlOP01&CtrlFunc10a)|(P1&CtrlOP01&CtrlFunc10b)|(P1&CtrlOP01&CtrlFunc10c)|(P1&CtrlOP01&CtrlFunc10e)|(P1&CtrlOP20)|(P1&CtrlOP21)|(P1&CtrlOP22)|(P1&CtrlOP23)|(P1&CtrlOP24)|(P1&CtrlOP25)|(P1&CtrlOP26)|(P1&CtrlOP30)|(P1&CtrlOP2b)|(P1&CtrlOP38)|(P1&CtrlOP00&CtrlFunc0b)|(P1&CtrlOP00&CtrlFunc0a)|(P1&CtrlOP00&CtrlFunc01)|(P1&CtrlOP1c&CtrlFunc20)|(P1&CtrlOP1c&CtrlFunc21)|(P1&CtrlOP11&CtrlFunc208)|(P1&CtrlOP10&CtrlFunc204)|(P1&CtrlOP11&CtrlFunc204)|(P1&CtrlOP1c&CtrlFunc00)|(P1&CtrlOP1c&CtrlFunc01)|(P1&CtrlOP1c&CtrlFunc04)|(P1&CtrlOP1c&CtrlFunc05)|(P1&CtrlOP28)|(P1&CtrlOP29)|(P1&CtrlOP2a)|(P1&CtrlOP2e);
assign CtrlALUOut=(P2&CtrlOP00&CtrlFunc20)|(P2&CtrlOP00&CtrlFunc22)|(P2&CtrlOP00&CtrlFunc21)|(P2&CtrlOP00&CtrlFunc23)|(P2&CtrlOP00&CtrlFunc24)|(P2&CtrlOP00&CtrlFunc25)|(P2&CtrlOP00&CtrlFunc26)|(P2&CtrlOP00&CtrlFunc27)|(P2&CtrlOP00&CtrlFunc2a)|(P2&CtrlOP00&CtrlFunc2b)|(P2&CtrlOP08)|(P2&CtrlOP09)|(P2&CtrlOP0a)|(P2&CtrlOP0b)|(P2&CtrlOP0c)|(P2&CtrlOP0d)|(P2&CtrlOP0e)|(P2&CtrlOP00&CtrlFunc04)|(P2&CtrlOP00&CtrlFunc06)|(P2&CtrlOP00&CtrlFunc07)|(P2&~nop&CtrlOP00&CtrlFunc00)|(P2&CtrlOP00&CtrlFunc02)|(P2&CtrlOP00&CtrlFunc03)|(P2&CtrlOP04)|(P2&CtrlOP05)|(P2&CtrlOP07)|(P2&CtrlOP06)|(P2&CtrlOP01)|(P2&CtrlOP01&CtrlFunc101)|(P2&CtrlOP01&CtrlFunc110)|(P2&CtrlOP01&CtrlFunc111)|(P2&CtrlOP20)|(P2&CtrlOP21)|(P2&CtrlOP22)|(P2&CtrlOP23)|(P2&CtrlOP24)|(P2&CtrlOP25)|(P2&CtrlOP26)|(P2&CtrlOP30)|(P2&CtrlOP2b)|(P2&CtrlOP38)|(P2&CtrlOP11&CtrlFunc208)|(P2&CtrlOP28)|(P2&CtrlOP29)|(P2&CtrlOP2a)|(P2&CtrlOP2e);
assign CtrlB=(P1&CtrlOP00&CtrlFunc20)|(P1&CtrlOP00&CtrlFunc22)|(P1&CtrlOP00&CtrlFunc21)|(P1&CtrlOP00&CtrlFunc23)|(P1&CtrlOP00&CtrlFunc24)|(P1&CtrlOP00&CtrlFunc25)|(P1&CtrlOP00&CtrlFunc26)|(P1&CtrlOP00&CtrlFunc27)|(P1&CtrlOP00&CtrlFunc2a)|(P1&CtrlOP00&CtrlFunc2b)|(P1&CtrlOP08)|(P1&CtrlOP09)|(P1&CtrlOP0a)|(P1&CtrlOP0b)|(P1&CtrlOP0c)|(P1&CtrlOP0d)|(P1&CtrlOP0e)|(P1&CtrlOP00&CtrlFunc04)|(P1&CtrlOP00&CtrlFunc06)|(P1&CtrlOP00&CtrlFunc07)|(P1&~nop&CtrlOP00&CtrlFunc00)|(P1&CtrlOP00&CtrlFunc02)|(P1&CtrlOP00&CtrlFunc03)|(P1&CtrlOP00&CtrlFunc18)|(P1&CtrlOP00&CtrlFunc19)|(P1&CtrlOP00&CtrlFunc1a)|(P1&CtrlOP00&CtrlFunc1b)|(P1&CtrlOP1c&CtrlFunc02)|(P1&CtrlOP04)|(P1&CtrlOP05)|(P1&CtrlOP07)|(P1&CtrlOP06)|(P1&CtrlOP01)|(P1&CtrlOP01&CtrlFunc101)|(P1&CtrlOP01&CtrlFunc110)|(P1&CtrlOP01&CtrlFunc111)|(P1&CtrlOP00&CtrlFunc30)|(P1&CtrlOP00&CtrlFunc31)|(P1&CtrlOP00&CtrlFunc32)|(P1&CtrlOP00&CtrlFunc33)|(P1&CtrlOP00&CtrlFunc34)|(P1&CtrlOP00&CtrlFunc36)|(P1&CtrlOP01&CtrlFunc108)|(P1&CtrlOP01&CtrlFunc109)|(P1&CtrlOP01&CtrlFunc10a)|(P1&CtrlOP01&CtrlFunc10b)|(P1&CtrlOP01&CtrlFunc10c)|(P1&CtrlOP01&CtrlFunc10e)|(P1&CtrlOP20)|(P1&CtrlOP21)|(P1&CtrlOP22)|(P3&CtrlOP22)|(P1&CtrlOP23)|(P1&CtrlOP24)|(P1&CtrlOP25)|(P1&CtrlOP26)|(P3&CtrlOP26)|(P1&CtrlOP30)|(P1&CtrlOP2b)|(P1&CtrlOP38)|(P1&CtrlOP00&CtrlFunc0b)|(P1&CtrlOP00&CtrlFunc0a)|(P1&CtrlOP1c&CtrlFunc00)|(P1&CtrlOP1c&CtrlFunc01)|(P1&CtrlOP1c&CtrlFunc04)|(P1&CtrlOP1c&CtrlFunc05)|(P1&CtrlOP28)|(P1&CtrlOP29)|(P1&CtrlOP2a)|(P1&CtrlOP2e);
assign CtrlCP0=(P2&CtrlOP10&CtrlFunc204);
assign CtrlCP0_ASID=(P1&CtrlOP10&CtrlFunc18)|(P1&CtrlOP00&CtrlFunc0c);
assign CtrlCP0_EPC=(P3&~lt&CtrlOP00&CtrlFunc30)|(P3&~lt&CtrlOP00&CtrlFunc31)|(P3&~lt&CtrlOP00&CtrlFunc32)|(P3&~lt&CtrlOP00&CtrlFunc33)|(P3&zero&CtrlOP00&CtrlFunc34)|(P3&~zero&CtrlOP00&CtrlFunc36)|(P3&~lt&CtrlOP01&CtrlFunc108)|(P3&~lt&CtrlOP01&CtrlFunc109)|(P3&lt&CtrlOP01&CtrlFunc10a)|(P3&lt&CtrlOP01&CtrlFunc10b)|(P3&zero&CtrlOP01&CtrlFunc10c)|(P3&~zero&CtrlOP01&CtrlFunc10e)|(P1&CtrlOP00&CtrlFunc0c)|(P1&CtrlOP00&CtrlFunc0d);
assign CtrlCP0_ExCode=(P3&~lt&CtrlOP00&CtrlFunc30)|(P3&~lt&CtrlOP00&CtrlFunc31)|(P3&~lt&CtrlOP00&CtrlFunc32)|(P3&~lt&CtrlOP00&CtrlFunc33)|(P3&zero&CtrlOP00&CtrlFunc34)|(P3&~zero&CtrlOP00&CtrlFunc36)|(P3&~lt&CtrlOP01&CtrlFunc108)|(P3&~lt&CtrlOP01&CtrlFunc109)|(P3&lt&CtrlOP01&CtrlFunc10a)|(P3&lt&CtrlOP01&CtrlFunc10b)|(P3&zero&CtrlOP01&CtrlFunc10c)|(P3&~zero&CtrlOP01&CtrlFunc10e)|(P1&CtrlOP00&CtrlFunc0c)|(P1&CtrlOP00&CtrlFunc0d);
assign CtrlCP1=(P2&CtrlOP11&CtrlFunc204);
assign CtrlConditionReg=(P2&CtrlOP04)|(P2&CtrlOP05)|(P2&CtrlOP07)|(P2&CtrlOP06)|(P2&CtrlOP01)|(P2&CtrlOP01&CtrlFunc101)|(P2&CtrlOP01&CtrlFunc110)|(P2&CtrlOP01&CtrlFunc111)|(P2&CtrlOP00&CtrlFunc30)|(P2&CtrlOP00&CtrlFunc31)|(P2&CtrlOP00&CtrlFunc32)|(P2&CtrlOP00&CtrlFunc33)|(P2&CtrlOP00&CtrlFunc34)|(P2&CtrlOP00&CtrlFunc36)|(P2&CtrlOP01&CtrlFunc108)|(P2&CtrlOP01&CtrlFunc109)|(P2&CtrlOP01&CtrlFunc10a)|(P2&CtrlOP01&CtrlFunc10b)|(P2&CtrlOP01&CtrlFunc10c)|(P2&CtrlOP01&CtrlFunc10e)|(P2&CtrlOP00&CtrlFunc0b)|(P2&CtrlOP00&CtrlFunc0a)|(P2&CtrlOP00&CtrlFunc01)|(P3&CtrlOP11&CtrlFunc208);
assign CtrlDMem=(P3&CtrlOP2b)|(P3&LLbit&CtrlOP38)|(P3&CtrlOP28)|(P3&CtrlOP29)|(P3&CtrlOP2a)|(P3&CtrlOP2e);
assign CtrlDR=(P3&CtrlOP20)|(P3&CtrlOP21)|(P3&CtrlOP22)|(P3&CtrlOP23)|(P3&CtrlOP24)|(P3&CtrlOP25)|(P3&CtrlOP26)|(P3&CtrlOP30)|(P1&CtrlOP2b)|(P1&CtrlOP38)|(P1&CtrlOP28)|(P2&CtrlOP29)|(P2&CtrlOP2a)|(P2&CtrlOP2e);
assign CtrlDR0=(P1&CtrlOP29)|(P1&CtrlOP2a)|(P1&CtrlOP2e);
assign CtrlGPR=(P4&~OV&CtrlOP00&CtrlFunc20)|(P4&~OV&CtrlOP00&CtrlFunc22)|(P4&CtrlOP00&CtrlFunc21)|(P4&CtrlOP00&CtrlFunc23)|(P4&CtrlOP00&CtrlFunc24)|(P4&CtrlOP00&CtrlFunc25)|(P4&CtrlOP00&CtrlFunc26)|(P4&CtrlOP00&CtrlFunc27)|(P4&CtrlOP00&CtrlFunc2a)|(P4&CtrlOP00&CtrlFunc2b)|(P4&~OV&CtrlOP08)|(P4&CtrlOP09)|(P4&CtrlOP0a)|(P4&CtrlOP0b)|(P4&CtrlOP0c)|(P4&CtrlOP0d)|(P4&CtrlOP0e)|(P4&CtrlOP00&CtrlFunc04)|(P4&CtrlOP00&CtrlFunc06)|(P4&CtrlOP00&CtrlFunc07)|(P4&~nop&CtrlOP00&CtrlFunc00)|(P4&CtrlOP00&CtrlFunc02)|(P4&CtrlOP00&CtrlFunc03)|(P4&CtrlOP1c&CtrlFunc02)|(P2&CtrlOP01&CtrlFunc110)|(P2&CtrlOP01&CtrlFunc111)|(P1&CtrlOP03)|(P1&CtrlOP00&CtrlFunc09)|(P4&CtrlOP20)|(P4&CtrlOP21)|(P4&CtrlOP22)|(P4&CtrlOP23)|(P4&CtrlOP24)|(P4&CtrlOP25)|(P4&CtrlOP26)|(P4&CtrlOP30)|(P4&CtrlOP38)|(P1&CtrlOP00&CtrlFunc10)|(P1&CtrlOP00&CtrlFunc12)|(P4&~zero&CtrlOP00&CtrlFunc0b)|(P4&zero&CtrlOP00&CtrlFunc0a)|(P4&fp&CtrlOP00&CtrlFunc01)|(P1&CtrlOP0f)|(P2&CtrlOP1c&CtrlFunc20)|(P2&CtrlOP1c&CtrlFunc21)|(P1&CtrlOP10&CtrlFunc200)|(P1&CtrlOP11&CtrlFunc200);
assign CtrlHi=(P2&CtrlOP00&CtrlFunc18)|(P2&CtrlOP00&CtrlFunc19)|(P2&CtrlOP00&CtrlFunc1a)|(P2&CtrlOP00&CtrlFunc1b)|(P1&CtrlOP00&CtrlFunc11)|(P2&CtrlOP1c&CtrlFunc00)|(P2&CtrlOP1c&CtrlFunc01)|(P2&CtrlOP1c&CtrlFunc04)|(P2&CtrlOP1c&CtrlFunc05);
assign CtrlIR=(P0);
assign CtrlLLbit=(P4&CtrlOP30);
assign CtrlLo=(P2&CtrlOP00&CtrlFunc18)|(P2&CtrlOP00&CtrlFunc19)|(P2&CtrlOP00&CtrlFunc1a)|(P2&CtrlOP00&CtrlFunc1b)|(P2&CtrlOP1c&CtrlFunc02)|(P1&CtrlOP00&CtrlFunc13)|(P2&CtrlOP1c&CtrlFunc00)|(P2&CtrlOP1c&CtrlFunc01)|(P2&CtrlOP1c&CtrlFunc04)|(P2&CtrlOP1c&CtrlFunc05);
assign CtrlMux10_1=(P0&CtrlOP10&CtrlFunc204)|(P0&CtrlOP11&CtrlFunc204);
assign CtrlMux10_2=(P0&CtrlOP00&CtrlFunc20)|(P0&CtrlOP00&CtrlFunc22)|(P0&CtrlOP00&CtrlFunc21)|(P0&CtrlOP00&CtrlFunc23)|(P0&CtrlOP00&CtrlFunc24)|(P0&CtrlOP00&CtrlFunc25)|(P0&CtrlOP00&CtrlFunc26)|(P0&CtrlOP00&CtrlFunc27)|(P0&CtrlOP00&CtrlFunc2a)|(P0&CtrlOP00&CtrlFunc2b)|(P0&CtrlOP08)|(P0&CtrlOP09)|(P0&CtrlOP0a)|(P0&CtrlOP0b)|(P0&CtrlOP0c)|(P0&CtrlOP0d)|(P0&CtrlOP0e)|(P0&CtrlOP00&CtrlFunc04)|(P0&CtrlOP00&CtrlFunc06)|(P0&CtrlOP00&CtrlFunc07)|(P0&CtrlOP00&CtrlFunc18)|(P0&CtrlOP00&CtrlFunc19)|(P0&CtrlOP00&CtrlFunc1a)|(P0&CtrlOP00&CtrlFunc1b)|(P0&CtrlOP1c&CtrlFunc02)|(P0&CtrlOP04)|(P0&CtrlOP05)|(P0&CtrlOP07)|(P0&CtrlOP06)|(P0&CtrlOP01)|(P0&CtrlOP01&CtrlFunc101)|(P0&CtrlOP01&CtrlFunc110)|(P0&CtrlOP01&CtrlFunc111)|(P0&CtrlOP00&CtrlFunc08)|(P0&CtrlOP00&CtrlFunc09)|(P0&CtrlOP00&CtrlFunc30)|(P0&CtrlOP00&CtrlFunc31)|(P0&CtrlOP00&CtrlFunc32)|(P0&CtrlOP00&CtrlFunc33)|(P0&CtrlOP00&CtrlFunc34)|(P0&CtrlOP00&CtrlFunc36)|(P0&CtrlOP01&CtrlFunc108)|(P0&CtrlOP01&CtrlFunc109)|(P0&CtrlOP01&CtrlFunc10a)|(P0&CtrlOP01&CtrlFunc10b)|(P0&CtrlOP01&CtrlFunc10c)|(P0&CtrlOP01&CtrlFunc10e)|(P0&CtrlOP20)|(P0&CtrlOP21)|(P0&CtrlOP22)|(P0&CtrlOP23)|(P0&CtrlOP24)|(P0&CtrlOP25)|(P0&CtrlOP26)|(P0&CtrlOP30)|(P0&CtrlOP2b)|(P0&CtrlOP38)|(P0&CtrlOP00&CtrlFunc11)|(P0&CtrlOP00&CtrlFunc13)|(P0&CtrlOP00&CtrlFunc0b)|(P0&CtrlOP00&CtrlFunc0a)|(P0&CtrlOP00&CtrlFunc01)|(P0&CtrlOP1c&CtrlFunc20)|(P0&CtrlOP1c&CtrlFunc21)|(P0&CtrlOP1c&CtrlFunc00)|(P0&CtrlOP1c&CtrlFunc01)|(P0&CtrlOP1c&CtrlFunc04)|(P0&CtrlOP1c&CtrlFunc05)|(P0&CtrlOP28)|(P0&CtrlOP29)|(P0&CtrlOP2a)|(P0&CtrlOP2e);
assign CtrlMux11_1=(P0&CtrlOP00&CtrlFunc20)|(P0&CtrlOP00&CtrlFunc22)|(P0&CtrlOP00&CtrlFunc21)|(P0&CtrlOP00&CtrlFunc23)|(P0&CtrlOP00&CtrlFunc24)|(P0&CtrlOP00&CtrlFunc25)|(P0&CtrlOP00&CtrlFunc26)|(P0&CtrlOP00&CtrlFunc27)|(P0&CtrlOP00&CtrlFunc2a)|(P0&CtrlOP00&CtrlFunc2b)|(P0&CtrlOP00&CtrlFunc04)|(P0&CtrlOP00&CtrlFunc06)|(P0&CtrlOP00&CtrlFunc07)|(P0&CtrlOP00&CtrlFunc00)|(P0&CtrlOP00&CtrlFunc02)|(P0&CtrlOP00&CtrlFunc03)|(P0&CtrlOP00&CtrlFunc18)|(P0&CtrlOP00&CtrlFunc19)|(P0&CtrlOP00&CtrlFunc1a)|(P0&CtrlOP00&CtrlFunc1b)|(P0&CtrlOP1c&CtrlFunc02)|(P0&CtrlOP04)|(P0&CtrlOP05)|(P0&CtrlOP07)|(P0&CtrlOP06)|(P0&CtrlOP01)|(P0&CtrlOP01&CtrlFunc101)|(P0&CtrlOP01&CtrlFunc110)|(P0&CtrlOP01&CtrlFunc111)|(P0&CtrlOP00&CtrlFunc30)|(P0&CtrlOP00&CtrlFunc31)|(P0&CtrlOP00&CtrlFunc32)|(P0&CtrlOP00&CtrlFunc33)|(P0&CtrlOP00&CtrlFunc34)|(P0&CtrlOP00&CtrlFunc36)|(P0&CtrlOP2b)|(P0&CtrlOP38)|(P0&CtrlOP00&CtrlFunc0b)|(P0&CtrlOP00&CtrlFunc0a)|(P0&CtrlOP1c&CtrlFunc00)|(P0&CtrlOP1c&CtrlFunc01)|(P0&CtrlOP1c&CtrlFunc04)|(P0&CtrlOP1c&CtrlFunc05)|(P0&CtrlOP28)|(P0&CtrlOP29)|(P0&CtrlOP2a)|(P0&CtrlOP2e)|(P2&CtrlOP22)|(P2&CtrlOP26);
assign CtrlMux12_1=(P3&CtrlOP00&CtrlFunc0b)|(P3&CtrlOP00&CtrlFunc0a)|(P3&CtrlOP00&CtrlFunc01);
assign CtrlMux12_10=(P0&CtrlOP03)|(P0&CtrlOP00&CtrlFunc09)|(P1&CtrlOP01&CtrlFunc110)|(P1&CtrlOP01&CtrlFunc111);
assign CtrlMux12_11=(P3&CtrlOP38);
assign CtrlMux12_2=(P3&CtrlOP00&CtrlFunc20)|(P3&CtrlOP00&CtrlFunc22)|(P3&CtrlOP00&CtrlFunc21)|(P3&CtrlOP00&CtrlFunc23)|(P3&CtrlOP00&CtrlFunc24)|(P3&CtrlOP00&CtrlFunc25)|(P3&CtrlOP00&CtrlFunc26)|(P3&CtrlOP00&CtrlFunc27)|(P3&CtrlOP00&CtrlFunc2a)|(P3&CtrlOP00&CtrlFunc2b)|(P3&CtrlOP08)|(P3&CtrlOP09)|(P3&CtrlOP0a)|(P3&CtrlOP0b)|(P3&CtrlOP0c)|(P3&CtrlOP0d)|(P3&CtrlOP0e)|(P3&CtrlOP00&CtrlFunc04)|(P3&CtrlOP00&CtrlFunc06)|(P3&CtrlOP00&CtrlFunc07)|(P3&~nop&CtrlOP00&CtrlFunc00)|(P3&CtrlOP00&CtrlFunc02)|(P3&CtrlOP00&CtrlFunc03);
assign CtrlMux12_3=(P0&CtrlOP10&CtrlFunc200);
assign CtrlMux12_4=(P0&CtrlOP11&CtrlFunc200);
assign CtrlMux12_5=(P1&CtrlOP1c&CtrlFunc20)|(P1&CtrlOP1c&CtrlFunc21);
assign CtrlMux12_6=(P0&CtrlOP00&CtrlFunc10);
assign CtrlMux12_7=(P0&CtrlOP0f);
assign CtrlMux12_8=(P0&CtrlOP00&CtrlFunc12)|(P3&CtrlOP1c&CtrlFunc02);
assign CtrlMux12_9=(P3&CtrlOP20)|(P3&CtrlOP21)|(P3&CtrlOP22)|(P3&CtrlOP23)|(P3&CtrlOP24)|(P3&CtrlOP25)|(P3&CtrlOP26)|(P3&CtrlOP30);
assign CtrlMux13_1=(P0&CtrlOP03)|(P1&CtrlOP01&CtrlFunc110)|(P1&CtrlOP01&CtrlFunc111);
assign CtrlMux13_2=(P0&CtrlOP00&CtrlFunc09)|(P0&CtrlOP00&CtrlFunc10)|(P0&CtrlOP00&CtrlFunc12)|(P1&CtrlOP1c&CtrlFunc20)|(P1&CtrlOP1c&CtrlFunc21)|(P3&CtrlOP00&CtrlFunc20)|(P3&CtrlOP00&CtrlFunc22)|(P3&CtrlOP00&CtrlFunc21)|(P3&CtrlOP00&CtrlFunc23)|(P3&CtrlOP00&CtrlFunc24)|(P3&CtrlOP00&CtrlFunc25)|(P3&CtrlOP00&CtrlFunc26)|(P3&CtrlOP00&CtrlFunc27)|(P3&CtrlOP00&CtrlFunc2a)|(P3&CtrlOP00&CtrlFunc2b)|(P3&CtrlOP00&CtrlFunc04)|(P3&CtrlOP00&CtrlFunc06)|(P3&CtrlOP00&CtrlFunc07)|(P3&~nop&CtrlOP00&CtrlFunc00)|(P3&CtrlOP00&CtrlFunc02)|(P3&CtrlOP00&CtrlFunc03)|(P3&CtrlOP1c&CtrlFunc02)|(P3&CtrlOP00&CtrlFunc0b)|(P3&CtrlOP00&CtrlFunc0a)|(P3&CtrlOP00&CtrlFunc01);
assign CtrlMux13_3=(P0&CtrlOP0f)|(P0&CtrlOP10&CtrlFunc200)|(P0&CtrlOP11&CtrlFunc200)|(P3&CtrlOP08)|(P3&CtrlOP09)|(P3&CtrlOP0a)|(P3&CtrlOP0b)|(P3&CtrlOP0c)|(P3&CtrlOP0d)|(P3&CtrlOP0e)|(P3&CtrlOP20)|(P3&CtrlOP21)|(P3&CtrlOP22)|(P3&CtrlOP23)|(P3&CtrlOP24)|(P3&CtrlOP25)|(P3&CtrlOP26)|(P3&CtrlOP30)|(P3&CtrlOP38);
assign CtrlMux14_1=(P0&CtrlOP00&CtrlFunc20)|(P0&CtrlOP00&CtrlFunc22)|(P0&CtrlOP00&CtrlFunc21)|(P0&CtrlOP00&CtrlFunc23)|(P0&CtrlOP00&CtrlFunc24)|(P0&CtrlOP00&CtrlFunc25)|(P0&CtrlOP00&CtrlFunc26)|(P0&CtrlOP00&CtrlFunc27)|(P0&CtrlOP00&CtrlFunc2a)|(P0&CtrlOP00&CtrlFunc2b)|(P0&CtrlOP08)|(P0&CtrlOP09)|(P0&CtrlOP0a)|(P0&CtrlOP0b)|(P0&CtrlOP0c)|(P0&CtrlOP0d)|(P0&CtrlOP0e)|(P0&CtrlOP00&CtrlFunc04)|(P0&CtrlOP00&CtrlFunc06)|(P0&CtrlOP00&CtrlFunc07)|(P0&CtrlOP00&CtrlFunc18)|(P0&CtrlOP00&CtrlFunc19)|(P0&CtrlOP00&CtrlFunc1a)|(P0&CtrlOP00&CtrlFunc1b)|(P0&CtrlOP1c&CtrlFunc02)|(P0&CtrlOP04)|(P0&CtrlOP05)|(P0&CtrlOP07)|(P0&CtrlOP06)|(P0&CtrlOP01)|(P0&CtrlOP01&CtrlFunc101)|(P0&CtrlOP01&CtrlFunc110)|(P0&CtrlOP01&CtrlFunc111)|(P0&CtrlOP00&CtrlFunc30)|(P0&CtrlOP00&CtrlFunc31)|(P0&CtrlOP00&CtrlFunc32)|(P0&CtrlOP00&CtrlFunc33)|(P0&CtrlOP00&CtrlFunc34)|(P0&CtrlOP00&CtrlFunc36)|(P0&CtrlOP01&CtrlFunc108)|(P0&CtrlOP01&CtrlFunc109)|(P0&CtrlOP01&CtrlFunc10a)|(P0&CtrlOP01&CtrlFunc10b)|(P0&CtrlOP01&CtrlFunc10c)|(P0&CtrlOP01&CtrlFunc10e)|(P0&CtrlOP20)|(P0&CtrlOP21)|(P0&CtrlOP22)|(P0&CtrlOP23)|(P0&CtrlOP24)|(P0&CtrlOP25)|(P0&CtrlOP26)|(P0&CtrlOP30)|(P0&CtrlOP2b)|(P0&CtrlOP38)|(P0&CtrlOP00&CtrlFunc0b)|(P0&CtrlOP00&CtrlFunc0a)|(P0&CtrlOP00&CtrlFunc01)|(P0&CtrlOP1c&CtrlFunc20)|(P0&CtrlOP1c&CtrlFunc21)|(P0&CtrlOP10&CtrlFunc204)|(P0&CtrlOP11&CtrlFunc204)|(P0&CtrlOP1c&CtrlFunc00)|(P0&CtrlOP1c&CtrlFunc01)|(P0&CtrlOP1c&CtrlFunc04)|(P0&CtrlOP1c&CtrlFunc05)|(P0&CtrlOP28)|(P0&CtrlOP29)|(P0&CtrlOP2a)|(P0&CtrlOP2e);
assign CtrlMux14_2=(P0&CtrlOP11&CtrlFunc208);
assign CtrlMux15_1=(P0&CtrlOP00&CtrlFunc20)|(P0&CtrlOP00&CtrlFunc22)|(P0&CtrlOP00&CtrlFunc21)|(P0&CtrlOP00&CtrlFunc23)|(P0&CtrlOP00&CtrlFunc24)|(P0&CtrlOP00&CtrlFunc25)|(P0&CtrlOP00&CtrlFunc26)|(P0&CtrlOP00&CtrlFunc27)|(P0&CtrlOP00&CtrlFunc2a)|(P0&CtrlOP00&CtrlFunc2b)|(P0&CtrlOP00&CtrlFunc04)|(P0&CtrlOP00&CtrlFunc06)|(P0&CtrlOP00&CtrlFunc07)|(P0&CtrlOP00&CtrlFunc00)|(P0&CtrlOP00&CtrlFunc02)|(P0&CtrlOP00&CtrlFunc03)|(P0&CtrlOP00&CtrlFunc18)|(P0&CtrlOP00&CtrlFunc19)|(P0&CtrlOP00&CtrlFunc1a)|(P0&CtrlOP00&CtrlFunc1b)|(P0&CtrlOP1c&CtrlFunc02)|(P0&CtrlOP04)|(P0&CtrlOP05)|(P0&CtrlOP07)|(P0&CtrlOP06)|(P0&CtrlOP01)|(P0&CtrlOP01&CtrlFunc101)|(P0&CtrlOP01&CtrlFunc110)|(P0&CtrlOP01&CtrlFunc111)|(P0&CtrlOP00&CtrlFunc30)|(P0&CtrlOP00&CtrlFunc31)|(P0&CtrlOP00&CtrlFunc32)|(P0&CtrlOP00&CtrlFunc33)|(P0&CtrlOP00&CtrlFunc34)|(P0&CtrlOP00&CtrlFunc36)|(P0&CtrlOP00&CtrlFunc0b)|(P0&CtrlOP00&CtrlFunc0a)|(P0&CtrlOP1c&CtrlFunc00)|(P0&CtrlOP1c&CtrlFunc01)|(P0&CtrlOP1c&CtrlFunc04)|(P0&CtrlOP1c&CtrlFunc05)|(P2&CtrlOP22)|(P2&CtrlOP26);
assign CtrlMux15_2=(P0&CtrlOP08)|(P0&CtrlOP09)|(P0&CtrlOP0a)|(P0&CtrlOP0b)|(P0&CtrlOP01&CtrlFunc108)|(P0&CtrlOP01&CtrlFunc109)|(P0&CtrlOP01&CtrlFunc10a)|(P0&CtrlOP01&CtrlFunc10b)|(P0&CtrlOP01&CtrlFunc10c)|(P0&CtrlOP01&CtrlFunc10e)|(P0&CtrlOP20)|(P0&CtrlOP21)|(P0&CtrlOP22)|(P0&CtrlOP23)|(P0&CtrlOP24)|(P0&CtrlOP25)|(P0&CtrlOP26)|(P0&CtrlOP30)|(P0&CtrlOP2b)|(P0&CtrlOP38)|(P0&CtrlOP28)|(P0&CtrlOP29)|(P0&CtrlOP2a)|(P0&CtrlOP2e);
assign CtrlMux15_3=(P0&CtrlOP0c)|(P0&CtrlOP0d)|(P0&CtrlOP0e);
assign CtrlMux16_1=(P1&CtrlOP00&CtrlFunc20)|(P1&CtrlOP00&CtrlFunc22)|(P1&CtrlOP00&CtrlFunc21)|(P1&CtrlOP00&CtrlFunc23)|(P1&CtrlOP00&CtrlFunc24)|(P1&CtrlOP00&CtrlFunc25)|(P1&CtrlOP00&CtrlFunc26)|(P1&CtrlOP00&CtrlFunc27)|(P1&CtrlOP00&CtrlFunc2a)|(P1&CtrlOP00&CtrlFunc2b)|(P1&CtrlOP08)|(P1&CtrlOP09)|(P1&CtrlOP0a)|(P1&CtrlOP0b)|(P1&CtrlOP0c)|(P1&CtrlOP0d)|(P1&CtrlOP0e)|(P1&CtrlOP20)|(P1&CtrlOP21)|(P1&CtrlOP22)|(P1&CtrlOP23)|(P1&CtrlOP24)|(P1&CtrlOP25)|(P1&CtrlOP26)|(P1&CtrlOP30)|(P1&CtrlOP2b)|(P1&CtrlOP38)|(P1&CtrlOP28)|(P1&CtrlOP29)|(P1&CtrlOP2a)|(P1&CtrlOP2e);
assign CtrlMux16_2=(P1&CtrlOP04)|(P1&CtrlOP05)|(P1&CtrlOP07)|(P1&CtrlOP06)|(P1&CtrlOP01)|(P1&CtrlOP01&CtrlFunc110)|(P1&CtrlOP01&CtrlFunc111)|(P1&CtrlOP11&CtrlFunc208);
assign CtrlMux16_3=(P1&CtrlOP01&CtrlFunc101);
assign CtrlMux17_1=(P1&CtrlOP00&CtrlFunc20)|(P1&CtrlOP00&CtrlFunc22)|(P1&CtrlOP00&CtrlFunc21)|(P1&CtrlOP00&CtrlFunc23)|(P1&CtrlOP00&CtrlFunc24)|(P1&CtrlOP00&CtrlFunc25)|(P1&CtrlOP00&CtrlFunc26)|(P1&CtrlOP00&CtrlFunc27)|(P1&CtrlOP00&CtrlFunc2a)|(P1&CtrlOP00&CtrlFunc2b)|(P1&CtrlOP08)|(P1&CtrlOP09)|(P1&CtrlOP0a)|(P1&CtrlOP0b)|(P1&CtrlOP0c)|(P1&CtrlOP0d)|(P1&CtrlOP0e)|(P1&CtrlOP20)|(P1&CtrlOP21)|(P1&CtrlOP22)|(P1&CtrlOP23)|(P1&CtrlOP24)|(P1&CtrlOP25)|(P1&CtrlOP26)|(P1&CtrlOP30)|(P1&CtrlOP2b)|(P1&CtrlOP38)|(P1&CtrlOP28)|(P1&CtrlOP29)|(P1&CtrlOP2a)|(P1&CtrlOP2e);
assign CtrlMux17_2=(P1&CtrlOP04)|(P1&CtrlOP05)|(P1&CtrlOP07)|(P1&CtrlOP06)|(P1&CtrlOP01)|(P1&CtrlOP01&CtrlFunc101)|(P1&CtrlOP01&CtrlFunc110)|(P1&CtrlOP01&CtrlFunc111)|(P1&CtrlOP11&CtrlFunc208);
assign CtrlMux18_1=(P1&CtrlOP00&CtrlFunc24)|(P1&CtrlOP0c);
assign CtrlMux18_2=(P1&CtrlOP00&CtrlFunc25)|(P1&CtrlOP0d);
assign CtrlMux18_3=(P1&CtrlOP00&CtrlFunc20)|(P1&CtrlOP00&CtrlFunc21)|(P1&CtrlOP08)|(P1&CtrlOP09);
assign CtrlMux18_4=(P1&CtrlOP00&CtrlFunc26)|(P1&CtrlOP0e);
assign CtrlMux18_5=(P1&CtrlOP00&CtrlFunc22)|(P1&CtrlOP00&CtrlFunc23);
assign CtrlMux18_6=(P1&CtrlOP00&CtrlFunc2b)|(P1&CtrlOP0b);
assign CtrlMux18_7=(P1&CtrlOP00&CtrlFunc27);
assign CtrlMux18_8=(P1&CtrlOP04)|(P1&CtrlOP05)|(P1&CtrlOP07)|(P1&CtrlOP06)|(P1&CtrlOP01)|(P1&CtrlOP01&CtrlFunc101)|(P1&CtrlOP01&CtrlFunc110)|(P1&CtrlOP01&CtrlFunc111)|(P1&CtrlOP20)|(P1&CtrlOP21)|(P1&CtrlOP22)|(P1&CtrlOP23)|(P1&CtrlOP24)|(P1&CtrlOP25)|(P1&CtrlOP26)|(P1&CtrlOP30)|(P1&CtrlOP2b)|(P1&CtrlOP38)|(P1&CtrlOP11&CtrlFunc208)|(P1&CtrlOP28)|(P1&CtrlOP29)|(P1&CtrlOP2a)|(P1&CtrlOP2e);
assign CtrlMux18_9=(P1&CtrlOP00&CtrlFunc2a)|(P1&CtrlOP0a);
assign CtrlMux19_1=(P1&CtrlOP00&CtrlFunc20)|(P1&CtrlOP00&CtrlFunc22)|(P1&CtrlOP00&CtrlFunc21)|(P1&CtrlOP00&CtrlFunc23)|(P1&CtrlOP00&CtrlFunc24)|(P1&CtrlOP00&CtrlFunc25)|(P1&CtrlOP00&CtrlFunc26)|(P1&CtrlOP00&CtrlFunc27)|(P1&CtrlOP00&CtrlFunc2a)|(P1&CtrlOP00&CtrlFunc2b)|(P1&CtrlOP08)|(P1&CtrlOP09)|(P1&CtrlOP0a)|(P1&CtrlOP0b)|(P1&CtrlOP0c)|(P1&CtrlOP0d)|(P1&CtrlOP0e)|(P1&CtrlOP04)|(P1&CtrlOP05)|(P1&CtrlOP07)|(P1&CtrlOP06)|(P1&CtrlOP01)|(P1&CtrlOP01&CtrlFunc101)|(P1&CtrlOP01&CtrlFunc110)|(P1&CtrlOP01&CtrlFunc111)|(P1&CtrlOP20)|(P1&CtrlOP21)|(P1&CtrlOP22)|(P1&CtrlOP23)|(P1&CtrlOP24)|(P1&CtrlOP25)|(P1&CtrlOP26)|(P1&CtrlOP30)|(P1&CtrlOP2b)|(P1&CtrlOP38)|(P1&CtrlOP11&CtrlFunc208)|(P1&CtrlOP28)|(P1&CtrlOP29)|(P1&CtrlOP2a)|(P1&CtrlOP2e);
assign CtrlMux19_2=(P1&CtrlOP00&CtrlFunc04)|(P1&CtrlOP00&CtrlFunc06)|(P1&CtrlOP00&CtrlFunc07)|(P1&~nop&CtrlOP00&CtrlFunc00)|(P1&CtrlOP00&CtrlFunc02)|(P1&CtrlOP00&CtrlFunc03);
assign CtrlMux1_1=(P0&CtrlOP02)|(P0&CtrlOP03);
assign CtrlMux1_2=(P3&CtrlOP04)|(P3&CtrlOP05)|(P3&CtrlOP07)|(P3&CtrlOP06)|(P3&CtrlOP01)|(P3&CtrlOP01&CtrlFunc101)|(P3&CtrlOP01&CtrlFunc110)|(P3&CtrlOP01&CtrlFunc111)|(P3&CtrlOP11&CtrlFunc208);
assign CtrlMux1_3=(P0&CtrlOP10&CtrlFunc18);
assign CtrlMux1_4=(P0&CtrlOP00&CtrlFunc0c)|(P0&CtrlOP00&CtrlFunc0d)|(P2&CtrlOP00&CtrlFunc30)|(P2&CtrlOP00&CtrlFunc31)|(P2&CtrlOP00&CtrlFunc32)|(P2&CtrlOP00&CtrlFunc33)|(P2&CtrlOP00&CtrlFunc34)|(P2&CtrlOP00&CtrlFunc36)|(P2&CtrlOP01&CtrlFunc108)|(P2&CtrlOP01&CtrlFunc109)|(P2&CtrlOP01&CtrlFunc10a)|(P2&CtrlOP01&CtrlFunc10b)|(P2&CtrlOP01&CtrlFunc10c)|(P2&CtrlOP01&CtrlFunc10e);
assign CtrlMux1_5=(P0&CtrlOP00&CtrlFunc08)|(P0&CtrlOP00&CtrlFunc09);
assign CtrlMux20_1=(P0&CtrlOP02)|(P0&CtrlOP03);
assign CtrlMux21_1=(P0&CtrlOP02)|(P0&CtrlOP03);
assign CtrlMux22_1=(P0&CtrlOP08)|(P0&CtrlOP09)|(P0&CtrlOP0a)|(P0&CtrlOP0b)|(P0&CtrlOP01&CtrlFunc108)|(P0&CtrlOP01&CtrlFunc109)|(P0&CtrlOP01&CtrlFunc10a)|(P0&CtrlOP01&CtrlFunc10b)|(P0&CtrlOP01&CtrlFunc10c)|(P0&CtrlOP01&CtrlFunc10e)|(P0&CtrlOP20)|(P0&CtrlOP21)|(P0&CtrlOP22)|(P0&CtrlOP23)|(P0&CtrlOP24)|(P0&CtrlOP25)|(P0&CtrlOP26)|(P0&CtrlOP30)|(P0&CtrlOP2b)|(P0&CtrlOP38)|(P0&CtrlOP28)|(P0&CtrlOP29)|(P0&CtrlOP2a)|(P0&CtrlOP2e);
assign CtrlMux23_1=(P0&CtrlOP0f);
assign CtrlMux24_1=(P0&CtrlOP0c)|(P0&CtrlOP0d)|(P0&CtrlOP0e);
assign CtrlMux25_1=(P0&CtrlOP11&CtrlFunc208)|(P1&CtrlOP04)|(P1&CtrlOP05)|(P1&CtrlOP07)|(P1&CtrlOP06)|(P1&CtrlOP01)|(P1&CtrlOP01&CtrlFunc101)|(P1&CtrlOP01&CtrlFunc110)|(P1&CtrlOP01&CtrlFunc111);
assign CtrlMux26_1=(P1&CtrlOP00&CtrlFunc0b)|(P1&CtrlOP00&CtrlFunc0a);
assign CtrlMux26_2=(P1&CtrlOP04)|(P1&CtrlOP05)|(P1&CtrlOP07)|(P1&CtrlOP06)|(P1&CtrlOP01)|(P1&CtrlOP01&CtrlFunc101)|(P1&CtrlOP01&CtrlFunc110)|(P1&CtrlOP01&CtrlFunc111)|(P1&CtrlOP00&CtrlFunc30)|(P1&CtrlOP00&CtrlFunc31)|(P1&CtrlOP00&CtrlFunc32)|(P1&CtrlOP00&CtrlFunc33)|(P1&CtrlOP00&CtrlFunc34)|(P1&CtrlOP00&CtrlFunc36)|(P1&CtrlOP01&CtrlFunc108)|(P1&CtrlOP01&CtrlFunc109)|(P1&CtrlOP01&CtrlFunc10a)|(P1&CtrlOP01&CtrlFunc10b)|(P1&CtrlOP01&CtrlFunc10c)|(P1&CtrlOP01&CtrlFunc10e);
assign CtrlMux27_1=(P1&CtrlOP04)|(P1&CtrlOP05)|(P1&CtrlOP07)|(P1&CtrlOP06)|(P1&CtrlOP01)|(P1&CtrlOP01&CtrlFunc101)|(P1&CtrlOP01&CtrlFunc110)|(P1&CtrlOP01&CtrlFunc111)|(P1&CtrlOP00&CtrlFunc30)|(P1&CtrlOP00&CtrlFunc31)|(P1&CtrlOP00&CtrlFunc32)|(P1&CtrlOP00&CtrlFunc33)|(P1&CtrlOP00&CtrlFunc34)|(P1&CtrlOP00&CtrlFunc36)|(P1&CtrlOP01&CtrlFunc108)|(P1&CtrlOP01&CtrlFunc109)|(P1&CtrlOP01&CtrlFunc10a)|(P1&CtrlOP01&CtrlFunc10b)|(P1&CtrlOP01&CtrlFunc10c)|(P1&CtrlOP01&CtrlFunc10e)|(P1&CtrlOP00&CtrlFunc0b)|(P1&CtrlOP00&CtrlFunc0a);
assign CtrlMux28_1=(P1&CtrlOP00&CtrlFunc31)|(P1&CtrlOP00&CtrlFunc33)|(P1&CtrlOP01&CtrlFunc109)|(P1&CtrlOP01&CtrlFunc10b);
assign CtrlMux28_2=(P1&CtrlOP04)|(P1&CtrlOP05)|(P1&CtrlOP07)|(P1&CtrlOP06)|(P1&CtrlOP01)|(P1&CtrlOP01&CtrlFunc101)|(P1&CtrlOP01&CtrlFunc110)|(P1&CtrlOP01&CtrlFunc111)|(P1&CtrlOP00&CtrlFunc30)|(P1&CtrlOP00&CtrlFunc32)|(P1&CtrlOP00&CtrlFunc34)|(P1&CtrlOP00&CtrlFunc36)|(P1&CtrlOP01&CtrlFunc108)|(P1&CtrlOP01&CtrlFunc10a)|(P1&CtrlOP01&CtrlFunc10c)|(P1&CtrlOP01&CtrlFunc10e)|(P1&CtrlOP00&CtrlFunc0b)|(P1&CtrlOP00&CtrlFunc0a);
assign CtrlMux29_1=(P1&CtrlOP1c&CtrlFunc20);
assign CtrlMux29_2=(P1&CtrlOP1c&CtrlFunc21);
assign CtrlMux2_1=((Reset|P4));
assign CtrlMux30_1=(P1&CtrlOP1c&CtrlFunc20)|(P1&CtrlOP1c&CtrlFunc21);
assign CtrlMux31_1=(P1&CtrlOP29)|(P1&CtrlOP2a)|(P1&CtrlOP2e)|(P2&CtrlOP20)|(P2&CtrlOP21)|(P2&CtrlOP22)|(P2&CtrlOP23)|(P2&CtrlOP24)|(P2&CtrlOP25)|(P2&CtrlOP26)|(P2&CtrlOP30);
assign CtrlMux31_2=(P0&CtrlOP2b)|(P0&CtrlOP38);
assign CtrlMux31_3=(P0&CtrlOP28);
assign CtrlMux32_1=(P0&CtrlOP29)|(P0&CtrlOP2a)|(P0&CtrlOP2e);
assign CtrlMux33_1=(P0&CtrlOP00&CtrlFunc11);
assign CtrlMux33_2=(P1&CtrlOP00&CtrlFunc18)|(P1&CtrlOP00&CtrlFunc19)|(P1&CtrlOP00&CtrlFunc1a)|(P1&CtrlOP00&CtrlFunc1b)|(P1&CtrlOP1c&CtrlFunc00)|(P1&CtrlOP1c&CtrlFunc01)|(P1&CtrlOP1c&CtrlFunc04)|(P1&CtrlOP1c&CtrlFunc05);
assign CtrlMux34_1=(P0&CtrlOP00&CtrlFunc13);
assign CtrlMux34_2=(P1&CtrlOP00&CtrlFunc18)|(P1&CtrlOP00&CtrlFunc19)|(P1&CtrlOP00&CtrlFunc1a)|(P1&CtrlOP00&CtrlFunc1b)|(P1&CtrlOP1c&CtrlFunc02)|(P1&CtrlOP1c&CtrlFunc00)|(P1&CtrlOP1c&CtrlFunc01)|(P1&CtrlOP1c&CtrlFunc04)|(P1&CtrlOP1c&CtrlFunc05);
assign CtrlMux35_1=(P3&CtrlOP30);
assign CtrlMux36_1=(P1&CtrlOP00&CtrlFunc18)|(P1&CtrlOP00&CtrlFunc19)|(P1&CtrlOP00&CtrlFunc1a)|(P1&CtrlOP00&CtrlFunc1b)|(P1&CtrlOP1c&CtrlFunc02)|(P1&CtrlOP1c&CtrlFunc00)|(P1&CtrlOP1c&CtrlFunc01)|(P1&CtrlOP1c&CtrlFunc04)|(P1&CtrlOP1c&CtrlFunc05);
assign CtrlMux37_1=(P1&CtrlOP00&CtrlFunc18)|(P1&CtrlOP00&CtrlFunc19)|(P1&CtrlOP00&CtrlFunc1a)|(P1&CtrlOP00&CtrlFunc1b)|(P1&CtrlOP1c&CtrlFunc02)|(P1&CtrlOP1c&CtrlFunc00)|(P1&CtrlOP1c&CtrlFunc01)|(P1&CtrlOP1c&CtrlFunc04)|(P1&CtrlOP1c&CtrlFunc05);
assign CtrlMux38_1=(P1&CtrlOP00&CtrlFunc18)|(P1&CtrlOP1c&CtrlFunc02);
assign CtrlMux38_2=(P1&CtrlOP00&CtrlFunc19);
assign CtrlMux38_3=(P1&CtrlOP00&CtrlFunc1a);
assign CtrlMux38_4=(P1&CtrlOP00&CtrlFunc1b);
assign CtrlMux38_5=(P1&CtrlOP1c&CtrlFunc00);
assign CtrlMux38_6=(P1&CtrlOP1c&CtrlFunc01);
assign CtrlMux38_7=(P1&CtrlOP1c&CtrlFunc04);
assign CtrlMux38_8=(P1&CtrlOP1c&CtrlFunc05);
assign CtrlMux39_1=(P1&CtrlOP1c&CtrlFunc00)|(P1&CtrlOP1c&CtrlFunc01)|(P1&CtrlOP1c&CtrlFunc04)|(P1&CtrlOP1c&CtrlFunc05);
assign CtrlMux3_1=((Reset|P4));
assign CtrlMux40_1=(P1&CtrlOP1c&CtrlFunc00)|(P1&CtrlOP1c&CtrlFunc01)|(P1&CtrlOP1c&CtrlFunc04)|(P1&CtrlOP1c&CtrlFunc05);
assign CtrlMux41_1=(P3&CtrlOP24);
assign CtrlMux41_10=(P2&CtrlOP2a);
assign CtrlMux41_11=(P2&CtrlOP38);
assign CtrlMux41_2=(P3&CtrlOP25);
assign CtrlMux41_3=(P3&CtrlOP26);
assign CtrlMux41_4=(P3&CtrlOP22);
assign CtrlMux41_5=(P3&CtrlOP23)|(P3&CtrlOP30);
assign CtrlMux41_6=(P3&CtrlOP20);
assign CtrlMux41_7=(P3&CtrlOP21);
assign CtrlMux41_8=(P2&CtrlOP29);
assign CtrlMux41_9=(P2&CtrlOP2e);
assign CtrlMux42_1=(P2&CtrlOP38)|(P2&CtrlOP29)|(P2&CtrlOP2a)|(P2&CtrlOP2e)|(P3&CtrlOP20)|(P3&CtrlOP21)|(P3&CtrlOP22)|(P3&CtrlOP23)|(P3&CtrlOP24)|(P3&CtrlOP25)|(P3&CtrlOP26)|(P3&CtrlOP30);
assign CtrlMux43_1=(P2&CtrlOP38)|(P2&CtrlOP29)|(P2&CtrlOP2a)|(P2&CtrlOP2e)|(P3&CtrlOP20)|(P3&CtrlOP21)|(P3&CtrlOP22)|(P3&CtrlOP23)|(P3&CtrlOP24)|(P3&CtrlOP25)|(P3&CtrlOP26)|(P3&CtrlOP30);
assign CtrlMux44_1=(P3&CtrlOP22)|(P3&CtrlOP26);
assign CtrlMux44_2=(P2&CtrlOP29)|(P2&CtrlOP2a)|(P2&CtrlOP2e);
assign CtrlMux45_1=(P1&CtrlOP00&CtrlFunc20)|(P1&CtrlOP00&CtrlFunc22)|(P1&CtrlOP08);
assign CtrlMux46_1=(P1&CtrlOP07)|(P1&CtrlOP06);
assign CtrlMux46_2=(P1&CtrlOP01)|(P1&CtrlOP01&CtrlFunc101)|(P1&CtrlOP01&CtrlFunc110)|(P1&CtrlOP01&CtrlFunc111)|(P1&CtrlOP00&CtrlFunc30)|(P1&CtrlOP00&CtrlFunc31)|(P1&CtrlOP00&CtrlFunc32)|(P1&CtrlOP00&CtrlFunc33)|(P1&CtrlOP01&CtrlFunc108)|(P1&CtrlOP01&CtrlFunc109)|(P1&CtrlOP01&CtrlFunc10a)|(P1&CtrlOP01&CtrlFunc10b);
assign CtrlMux46_3=(P1&CtrlOP04)|(P1&CtrlOP05)|(P1&CtrlOP00&CtrlFunc34)|(P1&CtrlOP00&CtrlFunc36)|(P1&CtrlOP01&CtrlFunc10c)|(P1&CtrlOP01&CtrlFunc10e)|(P1&CtrlOP00&CtrlFunc0b)|(P1&CtrlOP00&CtrlFunc0a);
assign CtrlMux46_4=(P1&CtrlOP00&CtrlFunc01)|(P2&CtrlOP11&CtrlFunc208);
assign CtrlMux47_1=(P0&CtrlOP00&CtrlFunc0c)|(P0&CtrlOP00&CtrlFunc0d)|(P2&CtrlOP00&CtrlFunc30)|(P2&CtrlOP00&CtrlFunc31)|(P2&CtrlOP00&CtrlFunc32)|(P2&CtrlOP00&CtrlFunc33)|(P2&CtrlOP00&CtrlFunc34)|(P2&CtrlOP00&CtrlFunc36)|(P2&CtrlOP01&CtrlFunc108)|(P2&CtrlOP01&CtrlFunc109)|(P2&CtrlOP01&CtrlFunc10a)|(P2&CtrlOP01&CtrlFunc10b)|(P2&CtrlOP01&CtrlFunc10c)|(P2&CtrlOP01&CtrlFunc10e);
assign CtrlMux48_1=(P1&CtrlOP00&CtrlFunc04)|(P1&CtrlOP00&CtrlFunc06)|(P1&CtrlOP00&CtrlFunc07)|(P1&~nop&CtrlOP00&CtrlFunc00)|(P1&CtrlOP00&CtrlFunc02)|(P1&CtrlOP00&CtrlFunc03);
assign CtrlMux49_1=(P1&CtrlOP00&CtrlFunc04)|(P1&~nop&CtrlOP00&CtrlFunc00);
assign CtrlMux49_2=(P1&CtrlOP00&CtrlFunc06)|(P1&CtrlOP00&CtrlFunc02);
assign CtrlMux49_3=(P1&CtrlOP00&CtrlFunc07)|(P1&CtrlOP00&CtrlFunc03);
assign CtrlMux4_1=(P1&CtrlOP28)|(P1&CtrlOP29)|(P1&CtrlOP2a)|(P1&CtrlOP2e)|(P2&CtrlOP20)|(P2&CtrlOP21)|(P2&CtrlOP22)|(P2&CtrlOP23)|(P2&CtrlOP24)|(P2&CtrlOP25)|(P2&CtrlOP26)|(P2&CtrlOP30)|(P2&CtrlOP2b)|(P2&CtrlOP38)|(P2&CtrlOP28)|(P2&CtrlOP29)|(P2&CtrlOP2a)|(P2&CtrlOP2e);
assign CtrlMux50_1=(P1&CtrlOP00&CtrlFunc04)|(P1&CtrlOP00&CtrlFunc06)|(P1&CtrlOP00&CtrlFunc07);
assign CtrlMux50_2=(P1&~nop&CtrlOP00&CtrlFunc00)|(P1&CtrlOP00&CtrlFunc02)|(P1&CtrlOP00&CtrlFunc03);
assign CtrlMux51_1=(P0&CtrlOP00&CtrlFunc0c);
assign CtrlMux51_2=(P0&CtrlOP10&CtrlFunc18);
assign CtrlMux52_1=(P0&CtrlOP00&CtrlFunc0c)|(P0&CtrlOP00&CtrlFunc0d)|(P2&CtrlOP00&CtrlFunc30)|(P2&CtrlOP00&CtrlFunc31)|(P2&CtrlOP00&CtrlFunc32)|(P2&CtrlOP00&CtrlFunc33)|(P2&CtrlOP00&CtrlFunc34)|(P2&CtrlOP00&CtrlFunc36)|(P2&CtrlOP01&CtrlFunc108)|(P2&CtrlOP01&CtrlFunc109)|(P2&CtrlOP01&CtrlFunc10a)|(P2&CtrlOP01&CtrlFunc10b)|(P2&CtrlOP01&CtrlFunc10c)|(P2&CtrlOP01&CtrlFunc10e);
assign CtrlMux53_1=(P0&CtrlOP00&CtrlFunc0c)|(P0&CtrlOP00&CtrlFunc0d);
assign CtrlMux53_2=(P2&CtrlOP00&CtrlFunc30)|(P2&CtrlOP00&CtrlFunc31)|(P2&CtrlOP00&CtrlFunc32)|(P2&CtrlOP00&CtrlFunc33)|(P2&CtrlOP00&CtrlFunc34)|(P2&CtrlOP00&CtrlFunc36)|(P2&CtrlOP01&CtrlFunc108)|(P2&CtrlOP01&CtrlFunc109)|(P2&CtrlOP01&CtrlFunc10a)|(P2&CtrlOP01&CtrlFunc10b)|(P2&CtrlOP01&CtrlFunc10c)|(P2&CtrlOP01&CtrlFunc10e);
assign CtrlMux54_1=(P0&CtrlOP10&CtrlFunc200);
assign CtrlMux55_1=(P1&CtrlOP10&CtrlFunc204);
assign CtrlMux56_1=(P1&CtrlOP10&CtrlFunc204);
assign CtrlMux57_1=(P1&CtrlOP00&CtrlFunc01)|(P2&CtrlOP11&CtrlFunc208);
assign CtrlMux58_1=(P0&CtrlOP11&CtrlFunc200);
assign CtrlMux59_1=(P1&CtrlOP00&CtrlFunc01)|(P2&CtrlOP11&CtrlFunc208);
assign CtrlMux5_1=(P1&CtrlOP28)|(P1&CtrlOP29)|(P1&CtrlOP2a)|(P1&CtrlOP2e)|(P2&CtrlOP20)|(P2&CtrlOP21)|(P2&CtrlOP22)|(P2&CtrlOP23)|(P2&CtrlOP24)|(P2&CtrlOP25)|(P2&CtrlOP26)|(P2&CtrlOP30);
assign CtrlMux60_1=(P1&CtrlOP11&CtrlFunc204);
assign CtrlMux61_1=(P1&CtrlOP11&CtrlFunc204);
assign CtrlMux64_1=(P4&CtrlOP00&CtrlFunc01)|(P4&CtrlOP11&CtrlFunc208);
assign CtrlMux65_1=(P4&CtrlOP07)|(P4&CtrlOP06);
assign CtrlMux68_1=(P0&CtrlOP00&CtrlFunc00);
assign CtrlMux69_1=(P3&CtrlOP38);
assign CtrlMux6_1=(P2&CtrlOP2b)|(P2&CtrlOP38)|(P2&CtrlOP28)|(P2&CtrlOP29)|(P2&CtrlOP2a)|(P2&CtrlOP2e);
assign CtrlMux70_1=(P3&CtrlOP00&CtrlFunc30)|(P3&CtrlOP00&CtrlFunc31)|(P3&CtrlOP00&CtrlFunc32)|(P3&CtrlOP00&CtrlFunc33)|(P3&CtrlOP01&CtrlFunc108)|(P3&CtrlOP01&CtrlFunc109)|(P3&CtrlOP01&CtrlFunc10a)|(P3&CtrlOP01&CtrlFunc10b)|(P4&CtrlOP01)|(P4&CtrlOP01&CtrlFunc101)|(P4&CtrlOP01&CtrlFunc110)|(P4&CtrlOP01&CtrlFunc111);
assign CtrlMux71_1=(P4&CtrlOP00&CtrlFunc20)|(P4&CtrlOP00&CtrlFunc22)|(P4&CtrlOP08);
assign CtrlMux72_1=(P3&CtrlOP00&CtrlFunc34)|(P3&CtrlOP00&CtrlFunc36)|(P3&CtrlOP01&CtrlFunc10c)|(P3&CtrlOP01&CtrlFunc10e)|(P4&CtrlOP04)|(P4&CtrlOP05)|(P4&CtrlOP00&CtrlFunc0b)|(P4&CtrlOP00&CtrlFunc0a);
assign CtrlMux7_1=(P2&CtrlOP2b)|(P2&CtrlOP28);
assign CtrlMux7_2=(P2&CtrlOP38)|(P2&CtrlOP29)|(P2&CtrlOP2a)|(P2&CtrlOP2e);
assign CtrlMux9_1=((Reset|P4));
assign CtrlOVReg=(P2&CtrlOP00&CtrlFunc20)|(P2&CtrlOP00&CtrlFunc22)|(P2&CtrlOP08);
assign CtrlPC=(P4&zero&CtrlOP04)|(P4&~zero&CtrlOP05)|(P4&gt&CtrlOP07)|(P4&~gt&CtrlOP06)|(P4&lt&CtrlOP01)|(P4&~lt&CtrlOP01&CtrlFunc101)|(P4&lt&CtrlOP01&CtrlFunc110)|(P4&~lt&CtrlOP01&CtrlFunc111)|(P1&CtrlOP02)|(P1&CtrlOP03)|(P1&CtrlOP00&CtrlFunc08)|(P1&CtrlOP00&CtrlFunc09)|(P3&~lt&CtrlOP00&CtrlFunc30)|(P3&~lt&CtrlOP00&CtrlFunc31)|(P3&~lt&CtrlOP00&CtrlFunc32)|(P3&~lt&CtrlOP00&CtrlFunc33)|(P3&zero&CtrlOP00&CtrlFunc34)|(P3&~zero&CtrlOP00&CtrlFunc36)|(P3&~lt&CtrlOP01&CtrlFunc108)|(P3&~lt&CtrlOP01&CtrlFunc109)|(P3&lt&CtrlOP01&CtrlFunc10a)|(P3&lt&CtrlOP01&CtrlFunc10b)|(P3&zero&CtrlOP01&CtrlFunc10c)|(P3&~zero&CtrlOP01&CtrlFunc10e)|(P4&fp&CtrlOP11&CtrlFunc208)|(P1&CtrlOP10&CtrlFunc18)|(P1&CtrlOP00&CtrlFunc0c)|(P1&CtrlOP00&CtrlFunc0d);
assign CtrlPCInc=(P0);
assign CtrlPIDReg=(P3&~lt&CtrlOP00&CtrlFunc30)|(P3&~lt&CtrlOP00&CtrlFunc31)|(P3&~lt&CtrlOP00&CtrlFunc32)|(P3&~lt&CtrlOP00&CtrlFunc33)|(P3&zero&CtrlOP00&CtrlFunc34)|(P3&~zero&CtrlOP00&CtrlFunc36)|(P3&~lt&CtrlOP01&CtrlFunc108)|(P3&~lt&CtrlOP01&CtrlFunc109)|(P3&lt&CtrlOP01&CtrlFunc10a)|(P3&lt&CtrlOP01&CtrlFunc10b)|(P3&zero&CtrlOP01&CtrlFunc10c)|(P3&~zero&CtrlOP01&CtrlFunc10e)|(P1&CtrlOP00&CtrlFunc0c)|(P1&CtrlOP00&CtrlFunc0d);
endmodule
