module CPU(clr,clk);
input clk,clr;
wire [5:0]CU_Func;
wire CtrlPCInc;
wire [31:0]PC_Out;
wire [31:0]IMem_Out;
wire CtrlIR;
wire [31:0]IR_Out;
wire CtrlRegs;
wire [31:0]Regs_Rdata1;
wire [31:0]Regs_Rdata2;
wire CtrlA;
wire [31:0]A_Out;
wire CtrlB;
wire [31:0]B_Out;
wire CtrlALUOut;
wire [31:0]ALUOut_Out;
wire [31:0]ALU_Out;
wire ALU_OV;
wire [31:0]CP0_ASID;
wire CtrlOVReg;
wire OVReg_Out;
CU_module CU(.clr(clr),.clk(clk),.Op(IR_Out[31:26]),.IRFunc(IR_Out[5:0]),.OV(OVReg_Out),.Func(CU_Func),.CtrlA(CtrlA),.CtrlALUOut(CtrlALUOut),.CtrlB(CtrlB),.CtrlIR(CtrlIR),.CtrlOVReg(CtrlOVReg),.CtrlPCInc(CtrlPCInc),.CtrlRegs(CtrlRegs));
PC_module PC(.clr(clr),.CtrlPCInc(CtrlPCInc),.Out(PC_Out));
IMemory_module IMem(.clr(clr),.RAddr(PC_Out),.ASID(CP0_ASID),.Out(IMem_Out));
IR_module IR(.clr(clr),.In(IMem_Out),.CtrlIR(CtrlIR),.Out(IR_Out));
Regs_module Regs(.clr(clr),.CtrlRegs(CtrlRegs),.RReg1(IR_Out[25:21]),.RReg2(IR_Out[20:16]),.WReg(IR_Out[15:11]),.WData(ALUOut_Out),.Rdata1(Regs_Rdata1),.Rdata2(Regs_Rdata2));
A_module A(.clr(clr),.CtrlA(CtrlA),.In(Regs_Rdata1),.Out(A_Out));
B_module B(.clr(clr),.CtrlB(CtrlB),.In(Regs_Rdata2),.Out(B_Out));
ALUOut_module ALUOut(.clr(clr),.CtrlALUOut(CtrlALUOut),.In(ALU_Out),.Out(ALUOut_Out));
ALU_module ALU(.A(A_Out),.B(B_Out),.Func(CU_Func),.Out(ALU_Out),.OV(ALU_OV));
CP0_module CP0(.clr(clr),.ASID(CP0_ASID));
OVReg_module OVReg(.clr(clr),.CtrlOVReg(CtrlOVReg),.In(ALU_OV),.Out(OVReg_Out));
endmodule
