module Initial_model(clr,clk,P0,P1,P2,P3,P4,Reset,Op,IRFunc,IRFunc1,IRFunc2,IR,nop,TrapAddr,CtrlFunc00,CtrlFunc01,CtrlFunc02,CtrlFunc03,CtrlFunc04,CtrlFunc05,CtrlFunc06,CtrlFunc07,CtrlFunc08,CtrlFunc09,CtrlFunc0a,CtrlFunc0b,CtrlFunc0c,CtrlFunc0d,CtrlFunc10,CtrlFunc101,CtrlFunc108,CtrlFunc109,CtrlFunc10a,CtrlFunc10b,CtrlFunc10c,CtrlFunc10e,CtrlFunc11,CtrlFunc110,CtrlFunc111,CtrlFunc12,CtrlFunc13,CtrlFunc18,CtrlFunc19,CtrlFunc1a,CtrlFunc1b,CtrlFunc20,CtrlFunc200,CtrlFunc204,CtrlFunc208,CtrlFunc21,CtrlFunc22,CtrlFunc23,CtrlFunc24,CtrlFunc25,CtrlFunc26,CtrlFunc27,CtrlFunc2a,CtrlFunc2b,CtrlFunc30,CtrlFunc31,CtrlFunc32,CtrlFunc33,CtrlFunc34,CtrlFunc36,CtrlOP00,CtrlOP01,CtrlOP02,CtrlOP03,CtrlOP04,CtrlOP05,CtrlOP06,CtrlOP07,CtrlOP08,CtrlOP09,CtrlOP0a,CtrlOP0b,CtrlOP0c,CtrlOP0d,CtrlOP0e,CtrlOP0f,CtrlOP10,CtrlOP11,CtrlOP1c,CtrlOP20,CtrlOP21,CtrlOP22,CtrlOP23,CtrlOP24,CtrlOP25,CtrlOP26,CtrlOP28,CtrlOP29,CtrlOP2a,CtrlOP2b,CtrlOP2e,CtrlOP30,CtrlOP38);
input clr,clk;
output P0;
output P1;
output P2;
output P3;
output P4;
output Reset;
input [5:0]Op;
input [5:0]IRFunc;
input [4:0]IRFunc1;
input [4:0]IRFunc2;
input [31:0]IR;
output nop;
output [31:0]TrapAddr;
output CtrlFunc00;
output CtrlFunc01;
output CtrlFunc02;
output CtrlFunc03;
output CtrlFunc04;
output CtrlFunc05;
output CtrlFunc06;
output CtrlFunc07;
output CtrlFunc08;
output CtrlFunc09;
output CtrlFunc0a;
output CtrlFunc0b;
output CtrlFunc0c;
output CtrlFunc0d;
output CtrlFunc10;
output CtrlFunc101;
output CtrlFunc108;
output CtrlFunc109;
output CtrlFunc10a;
output CtrlFunc10b;
output CtrlFunc10c;
output CtrlFunc10e;
output CtrlFunc11;
output CtrlFunc110;
output CtrlFunc111;
output CtrlFunc12;
output CtrlFunc13;
output CtrlFunc18;
output CtrlFunc19;
output CtrlFunc1a;
output CtrlFunc1b;
output CtrlFunc20;
output CtrlFunc200;
output CtrlFunc204;
output CtrlFunc208;
output CtrlFunc21;
output CtrlFunc22;
output CtrlFunc23;
output CtrlFunc24;
output CtrlFunc25;
output CtrlFunc26;
output CtrlFunc27;
output CtrlFunc2a;
output CtrlFunc2b;
output CtrlFunc30;
output CtrlFunc31;
output CtrlFunc32;
output CtrlFunc33;
output CtrlFunc34;
output CtrlFunc36;
output CtrlOP00;
output CtrlOP01;
output CtrlOP02;
output CtrlOP03;
output CtrlOP04;
output CtrlOP05;
output CtrlOP06;
output CtrlOP07;
output CtrlOP08;
output CtrlOP09;
output CtrlOP0a;
output CtrlOP0b;
output CtrlOP0c;
output CtrlOP0d;
output CtrlOP0e;
output CtrlOP0f;
output CtrlOP10;
output CtrlOP11;
output CtrlOP1c;
output CtrlOP20;
output CtrlOP21;
output CtrlOP22;
output CtrlOP23;
output CtrlOP24;
output CtrlOP25;
output CtrlOP26;
output CtrlOP28;
output CtrlOP29;
output CtrlOP2a;
output CtrlOP2b;
output CtrlOP2e;
output CtrlOP30;
output CtrlOP38;

wire [2:0]clkCounterOut;
Counter count(.clk(clk),.clr(clr),.dataout(clkCounterOut));
CP_generate clkgen(.dataIn(clkCounterOut),.Reset(Reset),.p0(P0),.p1(P1),.p2(P2),.p3(P3),.p4(P4));
assign CtrlFunc00=~IRFunc[5]&~IRFunc[4]&~IRFunc[3]&~IRFunc[2]&~IRFunc[1]&~IRFunc[0];
assign CtrlFunc01=~IRFunc[5]&~IRFunc[4]&~IRFunc[3]&~IRFunc[2]&~IRFunc[1]&IRFunc[0];
assign CtrlFunc02=~IRFunc[5]&~IRFunc[4]&~IRFunc[3]&~IRFunc[2]&IRFunc[1]&~IRFunc[0];
assign CtrlFunc03=~IRFunc[5]&~IRFunc[4]&~IRFunc[3]&~IRFunc[2]&IRFunc[1]&IRFunc[0];
assign CtrlFunc04=~IRFunc[5]&~IRFunc[4]&~IRFunc[3]&IRFunc[2]&~IRFunc[1]&~IRFunc[0];
assign CtrlFunc05=~IRFunc[5]&~IRFunc[4]&~IRFunc[3]&IRFunc[2]&~IRFunc[1]&IRFunc[0];
assign CtrlFunc06=~IRFunc[5]&~IRFunc[4]&~IRFunc[3]&IRFunc[2]&IRFunc[1]&~IRFunc[0];
assign CtrlFunc07=~IRFunc[5]&~IRFunc[4]&~IRFunc[3]&IRFunc[2]&IRFunc[1]&IRFunc[0];
assign CtrlFunc08=~IRFunc[5]&~IRFunc[4]&IRFunc[3]&~IRFunc[2]&~IRFunc[1]&~IRFunc[0];
assign CtrlFunc09=~IRFunc[5]&~IRFunc[4]&IRFunc[3]&~IRFunc[2]&~IRFunc[1]&IRFunc[0];
assign CtrlFunc0a=~IRFunc[5]&~IRFunc[4]&IRFunc[3]&~IRFunc[2]&IRFunc[1]&~IRFunc[0];
assign CtrlFunc0b=~IRFunc[5]&~IRFunc[4]&IRFunc[3]&~IRFunc[2]&IRFunc[1]&IRFunc[0];
assign CtrlFunc0c=~IRFunc[5]&~IRFunc[4]&IRFunc[3]&IRFunc[2]&~IRFunc[1]&~IRFunc[0];
assign CtrlFunc0d=~IRFunc[5]&~IRFunc[4]&IRFunc[3]&IRFunc[2]&~IRFunc[1]&IRFunc[0];
assign CtrlFunc10=~IRFunc[5]&IRFunc[4]&~IRFunc[3]&~IRFunc[2]&~IRFunc[1]&~IRFunc[0];
assign CtrlFunc101=~IRFunc1[4]&~IRFunc1[3]&~IRFunc1[2]&~IRFunc1[1]&IRFunc1[0];
assign CtrlFunc108=~IRFunc1[4]&IRFunc1[3]&~IRFunc1[2]&~IRFunc1[1]&~IRFunc1[0];
assign CtrlFunc109=~IRFunc1[4]&IRFunc1[3]&~IRFunc1[2]&~IRFunc1[1]&IRFunc1[0];
assign CtrlFunc10a=~IRFunc1[4]&IRFunc1[3]&~IRFunc1[2]&IRFunc1[1]&~IRFunc1[0];
assign CtrlFunc10b=~IRFunc1[4]&IRFunc1[3]&~IRFunc1[2]&IRFunc1[1]&IRFunc1[0];
assign CtrlFunc10c=~IRFunc1[4]&IRFunc1[3]&IRFunc1[2]&~IRFunc1[1]&~IRFunc1[0];
assign CtrlFunc10e=~IRFunc1[4]&IRFunc1[3]&IRFunc1[2]&IRFunc1[1]&~IRFunc1[0];
assign CtrlFunc11=~IRFunc[5]&IRFunc[4]&~IRFunc[3]&~IRFunc[2]&~IRFunc[1]&IRFunc[0];
assign CtrlFunc110=IRFunc1[4]&~IRFunc1[3]&~IRFunc1[2]&~IRFunc1[1]&~IRFunc1[0];
assign CtrlFunc111=IRFunc1[4]&~IRFunc1[3]&~IRFunc1[2]&~IRFunc1[1]&IRFunc1[0];
assign CtrlFunc12=~IRFunc[5]&IRFunc[4]&~IRFunc[3]&~IRFunc[2]&IRFunc[1]&~IRFunc[0];
assign CtrlFunc13=~IRFunc[5]&IRFunc[4]&~IRFunc[3]&~IRFunc[2]&IRFunc[1]&IRFunc[0];
assign CtrlFunc18=~IRFunc[5]&IRFunc[4]&IRFunc[3]&~IRFunc[2]&~IRFunc[1]&~IRFunc[0];
assign CtrlFunc19=~IRFunc[5]&IRFunc[4]&IRFunc[3]&~IRFunc[2]&~IRFunc[1]&IRFunc[0];
assign CtrlFunc1a=~IRFunc[5]&IRFunc[4]&IRFunc[3]&~IRFunc[2]&IRFunc[1]&~IRFunc[0];
assign CtrlFunc1b=~IRFunc[5]&IRFunc[4]&IRFunc[3]&~IRFunc[2]&IRFunc[1]&IRFunc[0];
assign CtrlFunc20=IRFunc[5]&~IRFunc[4]&~IRFunc[3]&~IRFunc[2]&~IRFunc[1]&~IRFunc[0];
assign CtrlFunc200=~IRFunc2[4]&~IRFunc2[3]&~IRFunc2[2]&~IRFunc2[1]&~IRFunc2[0];
assign CtrlFunc204=~IRFunc2[4]&~IRFunc2[3]&IRFunc2[2]&~IRFunc2[1]&~IRFunc2[0];
assign CtrlFunc208=~IRFunc2[4]&IRFunc2[3]&~IRFunc2[2]&~IRFunc2[1]&~IRFunc2[0];
assign CtrlFunc21=IRFunc[5]&~IRFunc[4]&~IRFunc[3]&~IRFunc[2]&~IRFunc[1]&IRFunc[0];
assign CtrlFunc22=IRFunc[5]&~IRFunc[4]&~IRFunc[3]&~IRFunc[2]&IRFunc[1]&~IRFunc[0];
assign CtrlFunc23=IRFunc[5]&~IRFunc[4]&~IRFunc[3]&~IRFunc[2]&IRFunc[1]&IRFunc[0];
assign CtrlFunc24=IRFunc[5]&~IRFunc[4]&~IRFunc[3]&IRFunc[2]&~IRFunc[1]&~IRFunc[0];
assign CtrlFunc25=IRFunc[5]&~IRFunc[4]&~IRFunc[3]&IRFunc[2]&~IRFunc[1]&IRFunc[0];
assign CtrlFunc26=IRFunc[5]&~IRFunc[4]&~IRFunc[3]&IRFunc[2]&IRFunc[1]&~IRFunc[0];
assign CtrlFunc27=IRFunc[5]&~IRFunc[4]&~IRFunc[3]&IRFunc[2]&IRFunc[1]&IRFunc[0];
assign CtrlFunc2a=IRFunc[5]&~IRFunc[4]&IRFunc[3]&~IRFunc[2]&IRFunc[1]&~IRFunc[0];
assign CtrlFunc2b=IRFunc[5]&~IRFunc[4]&IRFunc[3]&~IRFunc[2]&IRFunc[1]&IRFunc[0];
assign CtrlFunc30=IRFunc[5]&IRFunc[4]&~IRFunc[3]&~IRFunc[2]&~IRFunc[1]&~IRFunc[0];
assign CtrlFunc31=IRFunc[5]&IRFunc[4]&~IRFunc[3]&~IRFunc[2]&~IRFunc[1]&IRFunc[0];
assign CtrlFunc32=IRFunc[5]&IRFunc[4]&~IRFunc[3]&~IRFunc[2]&IRFunc[1]&~IRFunc[0];
assign CtrlFunc33=IRFunc[5]&IRFunc[4]&~IRFunc[3]&~IRFunc[2]&IRFunc[1]&IRFunc[0];
assign CtrlFunc34=IRFunc[5]&IRFunc[4]&~IRFunc[3]&IRFunc[2]&~IRFunc[1]&~IRFunc[0];
assign CtrlFunc36=IRFunc[5]&IRFunc[4]&~IRFunc[3]&IRFunc[2]&IRFunc[1]&~IRFunc[0];
assign CtrlOP00=~Op[5]&~Op[4]&~Op[3]&~Op[2]&~Op[1]&~Op[0];
assign CtrlOP01=~Op[5]&~Op[4]&~Op[3]&~Op[2]&~Op[1]&Op[0];
assign CtrlOP02=~Op[5]&~Op[4]&~Op[3]&~Op[2]&Op[1]&~Op[0];
assign CtrlOP03=~Op[5]&~Op[4]&~Op[3]&~Op[2]&Op[1]&Op[0];
assign CtrlOP04=~Op[5]&~Op[4]&~Op[3]&Op[2]&~Op[1]&~Op[0];
assign CtrlOP05=~Op[5]&~Op[4]&~Op[3]&Op[2]&~Op[1]&Op[0];
assign CtrlOP06=~Op[5]&~Op[4]&~Op[3]&Op[2]&Op[1]&~Op[0];
assign CtrlOP07=~Op[5]&~Op[4]&~Op[3]&Op[2]&Op[1]&Op[0];
assign CtrlOP08=~Op[5]&~Op[4]&Op[3]&~Op[2]&~Op[1]&~Op[0];
assign CtrlOP09=~Op[5]&~Op[4]&Op[3]&~Op[2]&~Op[1]&Op[0];
assign CtrlOP0a=~Op[5]&~Op[4]&Op[3]&~Op[2]&Op[1]&~Op[0];
assign CtrlOP0b=~Op[5]&~Op[4]&Op[3]&~Op[2]&Op[1]&Op[0];
assign CtrlOP0c=~Op[5]&~Op[4]&Op[3]&Op[2]&~Op[1]&~Op[0];
assign CtrlOP0d=~Op[5]&~Op[4]&Op[3]&Op[2]&~Op[1]&Op[0];
assign CtrlOP0e=~Op[5]&~Op[4]&Op[3]&Op[2]&Op[1]&~Op[0];
assign CtrlOP0f=~Op[5]&~Op[4]&Op[3]&Op[2]&Op[1]&Op[0];
assign CtrlOP10=~Op[5]&Op[4]&~Op[3]&~Op[2]&~Op[1]&~Op[0];
assign CtrlOP11=~Op[5]&Op[4]&~Op[3]&~Op[2]&~Op[1]&Op[0];
assign CtrlOP1c=~Op[5]&Op[4]&Op[3]&Op[2]&~Op[1]&~Op[0];
assign CtrlOP20=Op[5]&~Op[4]&~Op[3]&~Op[2]&~Op[1]&~Op[0];
assign CtrlOP21=Op[5]&~Op[4]&~Op[3]&~Op[2]&~Op[1]&Op[0];
assign CtrlOP22=Op[5]&~Op[4]&~Op[3]&~Op[2]&Op[1]&~Op[0];
assign CtrlOP23=Op[5]&~Op[4]&~Op[3]&~Op[2]&Op[1]&Op[0];
assign CtrlOP24=Op[5]&~Op[4]&~Op[3]&Op[2]&~Op[1]&~Op[0];
assign CtrlOP25=Op[5]&~Op[4]&~Op[3]&Op[2]&~Op[1]&Op[0];
assign CtrlOP26=Op[5]&~Op[4]&~Op[3]&Op[2]&Op[1]&~Op[0];
assign CtrlOP28=Op[5]&~Op[4]&Op[3]&~Op[2]&~Op[1]&~Op[0];
assign CtrlOP29=Op[5]&~Op[4]&Op[3]&~Op[2]&~Op[1]&Op[0];
assign CtrlOP2a=Op[5]&~Op[4]&Op[3]&~Op[2]&Op[1]&~Op[0];
assign CtrlOP2b=Op[5]&~Op[4]&Op[3]&~Op[2]&Op[1]&Op[0];
assign CtrlOP2e=Op[5]&~Op[4]&Op[3]&Op[2]&Op[1]&~Op[0];
assign CtrlOP30=Op[5]&Op[4]&~Op[3]&~Op[2]&~Op[1]&~Op[0];
assign CtrlOP38=Op[5]&Op[4]&Op[3]&~Op[2]&~Op[1]&~Op[0];
assign nop=~IR[31]&~IR[30]&~IR[29]&~IR[28]&~IR[27]&~IR[26]&~IR[25]&~IR[24]&~IR[23]&~IR[22]&~IR[21]&~IR[20]&~IR[19]&~IR[18]&~IR[17]&~IR[16]&~IR[15]&~IR[14]&~IR[13]&~IR[12]&~IR[11]&~IR[10]&~IR[9]&~IR[8]&~IR[7]&~IR[6]&~IR[5]&~IR[4]&~IR[3]&~IR[2]&~IR[1]&~IR[0];
assign TrapAddr=32'h80000200;
endmodule
