module mipsCPU(clr,clk);
input clk,clr;
wire CtrlMux1_1;
wire CtrlMux1_2;
wire CtrlMux1_3;
wire CtrlMux1_4;
wire CtrlMux1_5;
wire [31:0]Mux1_Out;
wire CtrlMux2_1;
wire [7:0]Mux2_Out;
wire CtrlMux3_1;
wire [31:0]Mux3_Out;
wire CtrlMux4_1;
wire [7:0]Mux4_Out;
wire CtrlMux5_1;
wire [31:0]Mux5_Out;
wire CtrlMux6_1;
wire [31:0]Mux6_Out;
wire CtrlMux7_1;
wire CtrlMux7_2;
wire [31:0]Mux7_Out;
wire CtrlMux9_1;
wire [31:0]Mux9_Out;
wire CtrlMux10_1;
wire CtrlMux10_2;
wire [4:0]Mux10_Out;
wire CtrlMux11_1;
wire [4:0]Mux11_Out;
wire CtrlMux12_1;
wire CtrlMux12_2;
wire CtrlMux12_3;
wire CtrlMux12_4;
wire CtrlMux12_5;
wire CtrlMux12_6;
wire CtrlMux12_7;
wire CtrlMux12_8;
wire CtrlMux12_9;
wire CtrlMux12_10;
wire CtrlMux12_11;
wire [31:0]Mux12_Out;
wire CtrlMux13_1;
wire CtrlMux13_2;
wire CtrlMux13_3;
wire [4:0]Mux13_Out;
wire CtrlMux14_1;
wire CtrlMux14_2;
wire [31:0]Mux14_Out;
wire CtrlMux15_1;
wire CtrlMux15_2;
wire CtrlMux15_3;
wire [31:0]Mux15_Out;
wire CtrlMux16_1;
wire CtrlMux16_2;
wire CtrlMux16_3;
wire [31:0]Mux16_Out;
wire CtrlMux17_1;
wire CtrlMux17_2;
wire [31:0]Mux17_Out;
wire CtrlMux18_1;
wire CtrlMux18_2;
wire CtrlMux18_3;
wire CtrlMux18_4;
wire CtrlMux18_5;
wire CtrlMux18_6;
wire CtrlMux18_7;
wire CtrlMux18_8;
wire CtrlMux18_9;
wire [5:0]Mux18_Out;
wire CtrlMux19_1;
wire CtrlMux19_2;
wire [31:0]Mux19_Out;
wire CtrlMux20_1;
wire [25:0]Mux20_Out;
wire CtrlMux21_1;
wire [3:0]Mux21_Out;
wire CtrlMux22_1;
wire [15:0]Mux22_Out;
wire CtrlMux23_1;
wire [15:0]Mux23_Out;
wire CtrlMux24_1;
wire [15:0]Mux24_Out;
wire CtrlMux25_1;
wire [15:0]Mux25_Out;
wire CtrlMux26_1;
wire CtrlMux26_2;
wire [31:0]Mux26_Out;
wire CtrlMux27_1;
wire [31:0]Mux27_Out;
wire CtrlMux28_1;
wire CtrlMux28_2;
wire [5:0]Mux28_Out;
wire CtrlMux29_1;
wire CtrlMux29_2;
wire [5:0]Mux29_Out;
wire CtrlMux30_1;
wire [31:0]Mux30_Out;
wire CtrlMux31_1;
wire CtrlMux31_2;
wire CtrlMux31_3;
wire [31:0]Mux31_Out;
wire CtrlMux32_1;
wire [31:0]Mux32_Out;
wire CtrlMux33_1;
wire CtrlMux33_2;
wire [31:0]Mux33_Out;
wire CtrlMux34_1;
wire CtrlMux34_2;
wire [31:0]Mux34_Out;
wire CtrlMux35_1;
wire Mux35_Out;
wire CtrlMux36_1;
wire [31:0]Mux36_Out;
wire CtrlMux37_1;
wire [31:0]Mux37_Out;
wire CtrlMux38_1;
wire CtrlMux38_2;
wire CtrlMux38_3;
wire CtrlMux38_4;
wire CtrlMux38_5;
wire CtrlMux38_6;
wire CtrlMux38_7;
wire CtrlMux38_8;
wire [5:0]Mux38_Out;
wire CtrlMux39_1;
wire [31:0]Mux39_Out;
wire CtrlMux40_1;
wire [31:0]Mux40_Out;
wire CtrlMux41_1;
wire CtrlMux41_2;
wire CtrlMux41_3;
wire CtrlMux41_4;
wire CtrlMux41_5;
wire CtrlMux41_6;
wire CtrlMux41_7;
wire CtrlMux41_8;
wire CtrlMux41_9;
wire CtrlMux41_10;
wire CtrlMux41_11;
wire [5:0]Mux41_Out;
wire CtrlMux42_1;
wire [1:0]Mux42_Out;
wire CtrlMux43_1;
wire [31:0]Mux43_Out;
wire CtrlMux44_1;
wire CtrlMux44_2;
wire [31:0]Mux44_Out;
wire CtrlMux45_1;
wire Mux45_Out;
wire CtrlMux46_1;
wire CtrlMux46_2;
wire CtrlMux46_3;
wire CtrlMux46_4;
wire Mux46_Out;
wire CtrlMux47_1;
wire [7:0]Mux47_Out;
wire CtrlMux48_1;
wire [31:0]Mux48_Out;
wire CtrlMux49_1;
wire CtrlMux49_2;
wire CtrlMux49_3;
wire [5:0]Mux49_Out;
wire CtrlMux50_1;
wire CtrlMux50_2;
wire [4:0]Mux50_Out;
wire CtrlMux51_1;
wire CtrlMux51_2;
wire [7:0]Mux51_Out;
wire CtrlMux52_1;
wire [31:0]Mux52_Out;
wire CtrlMux53_1;
wire CtrlMux53_2;
wire [4:0]Mux53_Out;
wire CtrlMux54_1;
wire [4:0]Mux54_Out;
wire CtrlMux55_1;
wire [31:0]Mux55_Out;
wire CtrlMux56_1;
wire [4:0]Mux56_Out;
wire CtrlMux57_1;
wire [2:0]Mux57_Out;
wire CtrlMux58_1;
wire [4:0]Mux58_Out;
wire CtrlMux59_1;
wire Mux59_Out;
wire CtrlMux60_1;
wire [31:0]Mux60_Out;
wire CtrlMux61_1;
wire [4:0]Mux61_Out;
wire CtrlMux64_1;
wire Mux64_Out;
wire CtrlMux65_1;
wire Mux65_Out;
wire CtrlMux68_1;
wire [31:0]Mux68_Out;
wire CtrlMux69_1;
wire Mux69_Out;
wire CtrlMux70_1;
wire Mux70_Out;
wire CtrlMux71_1;
wire Mux71_Out;
wire CtrlMux72_1;
wire Mux72_Out;
wire [31:0]CU_TrapAddr;
wire CtrlPC;
wire CtrlPCInc;
wire [31:0]PC_CIA;
wire [31:0]PC_Out;
wire [31:0]IMem_Out;
wire CtrlDMem;
wire [31:0]DMem_Out;
wire CtrlIR;
wire [31:0]IR_Out;
wire CtrlGPR;
wire [31:0]GPR_Rdata1;
wire [31:0]GPR_Rdata2;
wire CtrlA;
wire [31:0]A_Out;
wire CtrlB;
wire [31:0]B_Out;
wire CtrlALUOut;
wire [31:0]ALUOut_Out;
wire [31:0]ALU_Out;
wire ALU_OV;
wire [31:0]SU_Out;
wire CMPU_zero;
wire CMPU_lt;
wire CMPU_gt;
wire [31:0]IMMEXT_Out;
wire [31:0]IMMSEXT_Out;
wire [31:0]LIMMEXT_Out;
wire [31:0]ADDREXT_Out;
wire [31:0]SEXT_Out;
wire [31:0]CountUnit_Out;
wire CtrlDR;
wire [31:0]DR_Out;
wire CtrlDR0;
wire [31:0]DR0_Out;
wire CtrlLLbit;
wire LLbit_Out;
wire CtrlPIDReg;
wire [7:0]PIDReg_Out;
wire CtrlHi;
wire [31:0]Hi_Out;
wire CtrlLo;
wire [31:0]Lo_Out;
wire [31:0]MDU_lo;
wire [31:0]MDU_hi;
wire [31:0]MemDataSel_Out;
wire CtrlCP0_EPC;
wire CtrlCP0_ASID;
wire CtrlCP0_ExCode;
wire CtrlCP0;
wire [31:0]CP0_Rdata;
wire [31:0]CP0_EPC;
wire [7:0]CP0_ASID;
wire CtrlCP1;
wire CP1_fp;
wire [31:0]CP1_Rdata;
wire CtrlOVReg;
wire OVReg_Out;
wire CtrlConditionReg;
wire ConditionReg_Out;
CU_module CU(.clr(clr),.clk(clk),.Op(IR_Out[31:26]),.IRFunc(IR_Out[5:0]),.IRFunc1(IR_Out[20:16]),.IRFunc2(IR_Out[25:21]),.zero(Mux72_Out),.OV(Mux71_Out),.lt(Mux70_Out),.gt(Mux65_Out),.LLbit(Mux69_Out),.fp(Mux64_Out),.IR(Mux68_Out),.TrapAddr(CU_TrapAddr),.CtrlA(CtrlA),.CtrlALUOut(CtrlALUOut),.CtrlB(CtrlB),.CtrlCP0(CtrlCP0),.CtrlCP0_ASID(CtrlCP0_ASID),.CtrlCP0_EPC(CtrlCP0_EPC),.CtrlCP0_ExCode(CtrlCP0_ExCode),.CtrlCP1(CtrlCP1),.CtrlConditionReg(CtrlConditionReg),.CtrlDMem(CtrlDMem),.CtrlDR(CtrlDR),.CtrlDR0(CtrlDR0),.CtrlGPR(CtrlGPR),.CtrlHi(CtrlHi),.CtrlIR(CtrlIR),.CtrlLLbit(CtrlLLbit),.CtrlLo(CtrlLo),.CtrlOVReg(CtrlOVReg),.CtrlPC(CtrlPC),.CtrlPCInc(CtrlPCInc),.CtrlPIDReg(CtrlPIDReg),.CtrlMux1_1(CtrlMux1_1),.CtrlMux1_2(CtrlMux1_2),.CtrlMux1_3(CtrlMux1_3),.CtrlMux1_4(CtrlMux1_4),.CtrlMux1_5(CtrlMux1_5),.CtrlMux2_1(CtrlMux2_1),.CtrlMux3_1(CtrlMux3_1),.CtrlMux4_1(CtrlMux4_1),.CtrlMux5_1(CtrlMux5_1),.CtrlMux6_1(CtrlMux6_1),.CtrlMux7_1(CtrlMux7_1),.CtrlMux7_2(CtrlMux7_2),.CtrlMux9_1(CtrlMux9_1),.CtrlMux10_1(CtrlMux10_1),.CtrlMux10_2(CtrlMux10_2),.CtrlMux11_1(CtrlMux11_1),.CtrlMux12_1(CtrlMux12_1),.CtrlMux12_2(CtrlMux12_2),.CtrlMux12_3(CtrlMux12_3),.CtrlMux12_4(CtrlMux12_4),.CtrlMux12_5(CtrlMux12_5),.CtrlMux12_6(CtrlMux12_6),.CtrlMux12_7(CtrlMux12_7),.CtrlMux12_8(CtrlMux12_8),.CtrlMux12_9(CtrlMux12_9),.CtrlMux12_10(CtrlMux12_10),.CtrlMux12_11(CtrlMux12_11),.CtrlMux13_1(CtrlMux13_1),.CtrlMux13_2(CtrlMux13_2),.CtrlMux13_3(CtrlMux13_3),.CtrlMux14_1(CtrlMux14_1),.CtrlMux14_2(CtrlMux14_2),.CtrlMux15_1(CtrlMux15_1),.CtrlMux15_2(CtrlMux15_2),.CtrlMux15_3(CtrlMux15_3),.CtrlMux16_1(CtrlMux16_1),.CtrlMux16_2(CtrlMux16_2),.CtrlMux16_3(CtrlMux16_3),.CtrlMux17_1(CtrlMux17_1),.CtrlMux17_2(CtrlMux17_2),.CtrlMux18_1(CtrlMux18_1),.CtrlMux18_2(CtrlMux18_2),.CtrlMux18_3(CtrlMux18_3),.CtrlMux18_4(CtrlMux18_4),.CtrlMux18_5(CtrlMux18_5),.CtrlMux18_6(CtrlMux18_6),.CtrlMux18_7(CtrlMux18_7),.CtrlMux18_8(CtrlMux18_8),.CtrlMux18_9(CtrlMux18_9),.CtrlMux19_1(CtrlMux19_1),.CtrlMux19_2(CtrlMux19_2),.CtrlMux20_1(CtrlMux20_1),.CtrlMux21_1(CtrlMux21_1),.CtrlMux22_1(CtrlMux22_1),.CtrlMux23_1(CtrlMux23_1),.CtrlMux24_1(CtrlMux24_1),.CtrlMux25_1(CtrlMux25_1),.CtrlMux26_1(CtrlMux26_1),.CtrlMux26_2(CtrlMux26_2),.CtrlMux27_1(CtrlMux27_1),.CtrlMux28_1(CtrlMux28_1),.CtrlMux28_2(CtrlMux28_2),.CtrlMux29_1(CtrlMux29_1),.CtrlMux29_2(CtrlMux29_2),.CtrlMux30_1(CtrlMux30_1),.CtrlMux31_1(CtrlMux31_1),.CtrlMux31_2(CtrlMux31_2),.CtrlMux31_3(CtrlMux31_3),.CtrlMux32_1(CtrlMux32_1),.CtrlMux33_1(CtrlMux33_1),.CtrlMux33_2(CtrlMux33_2),.CtrlMux34_1(CtrlMux34_1),.CtrlMux34_2(CtrlMux34_2),.CtrlMux35_1(CtrlMux35_1),.CtrlMux36_1(CtrlMux36_1),.CtrlMux37_1(CtrlMux37_1),.CtrlMux38_1(CtrlMux38_1),.CtrlMux38_2(CtrlMux38_2),.CtrlMux38_3(CtrlMux38_3),.CtrlMux38_4(CtrlMux38_4),.CtrlMux38_5(CtrlMux38_5),.CtrlMux38_6(CtrlMux38_6),.CtrlMux38_7(CtrlMux38_7),.CtrlMux38_8(CtrlMux38_8),.CtrlMux39_1(CtrlMux39_1),.CtrlMux40_1(CtrlMux40_1),.CtrlMux41_1(CtrlMux41_1),.CtrlMux41_2(CtrlMux41_2),.CtrlMux41_3(CtrlMux41_3),.CtrlMux41_4(CtrlMux41_4),.CtrlMux41_5(CtrlMux41_5),.CtrlMux41_6(CtrlMux41_6),.CtrlMux41_7(CtrlMux41_7),.CtrlMux41_8(CtrlMux41_8),.CtrlMux41_9(CtrlMux41_9),.CtrlMux41_10(CtrlMux41_10),.CtrlMux41_11(CtrlMux41_11),.CtrlMux42_1(CtrlMux42_1),.CtrlMux43_1(CtrlMux43_1),.CtrlMux44_1(CtrlMux44_1),.CtrlMux44_2(CtrlMux44_2),.CtrlMux45_1(CtrlMux45_1),.CtrlMux46_1(CtrlMux46_1),.CtrlMux46_2(CtrlMux46_2),.CtrlMux46_3(CtrlMux46_3),.CtrlMux46_4(CtrlMux46_4),.CtrlMux47_1(CtrlMux47_1),.CtrlMux48_1(CtrlMux48_1),.CtrlMux49_1(CtrlMux49_1),.CtrlMux49_2(CtrlMux49_2),.CtrlMux49_3(CtrlMux49_3),.CtrlMux50_1(CtrlMux50_1),.CtrlMux50_2(CtrlMux50_2),.CtrlMux51_1(CtrlMux51_1),.CtrlMux51_2(CtrlMux51_2),.CtrlMux52_1(CtrlMux52_1),.CtrlMux53_1(CtrlMux53_1),.CtrlMux53_2(CtrlMux53_2),.CtrlMux54_1(CtrlMux54_1),.CtrlMux55_1(CtrlMux55_1),.CtrlMux56_1(CtrlMux56_1),.CtrlMux57_1(CtrlMux57_1),.CtrlMux58_1(CtrlMux58_1),.CtrlMux59_1(CtrlMux59_1),.CtrlMux60_1(CtrlMux60_1),.CtrlMux61_1(CtrlMux61_1),.CtrlMux64_1(CtrlMux64_1),.CtrlMux65_1(CtrlMux65_1),.CtrlMux68_1(CtrlMux68_1),.CtrlMux69_1(CtrlMux69_1),.CtrlMux70_1(CtrlMux70_1),.CtrlMux71_1(CtrlMux71_1),.CtrlMux72_1(CtrlMux72_1));
PC_module PC(.clr(clr),.CtrlPC(CtrlPC),.CtrlPCInc(CtrlPCInc),.In(Mux1_Out),.CIA(PC_CIA),.Out(PC_Out));
IMemory_module IMem(.clr(clr),.CtrlIMem(1'b0),.RAddr(Mux3_Out),.ASID(Mux2_Out),.Out(IMem_Out));
DMemory_module DMem(.clr(clr),.CtrlDMem(CtrlDMem),.WData(Mux7_Out),.WAddr(Mux6_Out),.RAddr(Mux5_Out),.ASID(Mux4_Out),.Out(DMem_Out));
IR_module IR(.clr(clr),.In(Mux9_Out),.CtrlIR(CtrlIR),.Out(IR_Out));
GPR_module GPR(.clr(clr),.CtrlGPR(CtrlGPR),.RReg1(Mux10_Out),.RReg2(Mux11_Out),.WReg(Mux13_Out),.WData(Mux12_Out),.Rdata1(GPR_Rdata1),.Rdata2(GPR_Rdata2));
A_module A(.clr(clr),.CtrlA(CtrlA),.In(Mux14_Out),.Out(A_Out));
B_module B(.clr(clr),.CtrlB(CtrlB),.In(Mux15_Out),.Out(B_Out));
ALUOut_module ALUOut(.clr(clr),.CtrlALUOut(CtrlALUOut),.In(Mux19_Out),.Out(ALUOut_Out));
ALU_module ALU(.A(Mux16_Out),.B(Mux17_Out),.Func(Mux18_Out),.Out(ALU_Out),.OV(ALU_OV));
Shift_unit SU(.Data(Mux48_Out),.Shamt(Mux50_Out),.Func(Mux49_Out),.Out(SU_Out));
CMPU_module CMPU(.A(Mux26_Out),.B(Mux27_Out),.Func(Mux28_Out),.zero(CMPU_zero),.lt(CMPU_lt),.gt(CMPU_gt));
IMMEXT_module IMMEXT(.In(Mux22_Out),.Out(IMMEXT_Out));
IMMSEXT_module IMMSEXT(.In(Mux23_Out),.Out(IMMSEXT_Out));
LIMMEXT_module LIMMEXT(.In(Mux24_Out),.Out(LIMMEXT_Out));
ADDREXT_module ADDREXT(.In(Mux20_Out),.PCpart(Mux21_Out),.Out(ADDREXT_Out));
SEXT_module SEXT(.In(Mux25_Out),.Out(SEXT_Out));
CountUnit_module CountUnit(.In(Mux30_Out),.Func(Mux29_Out),.Out(CountUnit_Out));
DR_module DR(.clr(clr),.CtrlDR(CtrlDR),.In(Mux31_Out),.Out(DR_Out));
DR0_module DR0(.clr(clr),.CtrlDR0(CtrlDR0),.In(Mux32_Out),.Out(DR0_Out));
LLbit_module LLbit(.clr(clr),.CtrlLLbit(CtrlLLbit),.In(Mux35_Out),.Out(LLbit_Out));
PIDReg_module PIDReg(.clr(clr),.CtrlPIDReg(CtrlPIDReg),.In(Mux47_Out),.Out(PIDReg_Out));
Hi_module Hi(.clr(clr),.CtrlHi(CtrlHi),.In(Mux33_Out),.Out(Hi_Out));
Lo_module Lo(.clr(clr),.CtrlLo(CtrlLo),.In(Mux34_Out),.Out(Lo_Out));
MDU_module MDU(.Lo(Mux40_Out),.Hi(Mux39_Out),.A(Mux36_Out),.B(Mux37_Out),.Func(Mux38_Out),.lo(MDU_lo),.hi(MDU_hi));
MemDataSel_module MemDataSel(.In(Mux43_Out),.Func(Mux41_Out),.Addr(Mux42_Out),.GPRIn(Mux44_Out),.Out(MemDataSel_Out));
CP0_module CP0(.clr(clr),.WReg(Mux56_Out),.Wdata(Mux55_Out),.RReg(Mux54_Out),.ExCodeIn(Mux53_Out),.EPCIn(Mux52_Out),.ASIDIn(Mux51_Out),.CtrlCP0_EPC(CtrlCP0_EPC),.CtrlCP0_ASID(CtrlCP0_ASID),.CtrlCP0_ExCode(CtrlCP0_ExCode),.CtrlCP0(CtrlCP0),.Rdata(CP0_Rdata),.EPC(CP0_EPC),.ASID(CP0_ASID));
CP1_module CP1(.clr(clr),.WReg(Mux61_Out),.Wdata(Mux60_Out),.RReg(Mux58_Out),.tf(Mux59_Out),.cc(Mux57_Out),.CtrlCP1(CtrlCP1),.fp(CP1_fp),.Rdata(CP1_Rdata));
OVReg_module OVReg(.clr(clr),.CtrlOVReg(CtrlOVReg),.In(Mux45_Out),.Out(OVReg_Out));
ConditionReg_module ConditionReg(.clr(clr),.CtrlConditionReg(CtrlConditionReg),.In(Mux46_Out),.Out(ConditionReg_Out));
Mux5_32module Mux1(.Mux_1(ADDREXT_Out),.SelMux_1(CtrlMux1_1),.Mux_2(ALUOut_Out),.SelMux_2(CtrlMux1_2),.Mux_3(CP0_EPC),.SelMux_3(CtrlMux1_3),.Mux_4(CU_TrapAddr),.SelMux_4(CtrlMux1_4),.Mux_5(GPR_Rdata1),.SelMux_5(CtrlMux1_5),.Out(Mux1_Out));
Mux1_8module Mux2(.Mux_1(CP0_ASID),.SelMux_1(CtrlMux2_1),.Out(Mux2_Out));
Mux1_32module Mux3(.Mux_1(PC_Out),.SelMux_1(CtrlMux3_1),.Out(Mux3_Out));
Mux1_8module Mux4(.Mux_1(CP0_ASID),.SelMux_1(CtrlMux4_1),.Out(Mux4_Out));
Mux1_32module Mux5(.Mux_1(ALUOut_Out),.SelMux_1(CtrlMux5_1),.Out(Mux5_Out));
Mux1_32module Mux6(.Mux_1(ALUOut_Out),.SelMux_1(CtrlMux6_1),.Out(Mux6_Out));
Mux2_32module Mux7(.Mux_1(DR_Out),.SelMux_1(CtrlMux7_1),.Mux_2(MemDataSel_Out),.SelMux_2(CtrlMux7_2),.Out(Mux7_Out));
Mux1_32module Mux9(.Mux_1(IMem_Out),.SelMux_1(CtrlMux9_1),.Out(Mux9_Out));
Mux2_5module Mux10(.Mux_1(IR_Out[20:16]),.SelMux_1(CtrlMux10_1),.Mux_2(IR_Out[25:21]),.SelMux_2(CtrlMux10_2),.Out(Mux10_Out));
Mux1_5module Mux11(.Mux_1(IR_Out[20:16]),.SelMux_1(CtrlMux11_1),.Out(Mux11_Out));
Mux11_32module Mux12(.Mux_1(A_Out),.SelMux_1(CtrlMux12_1),.Mux_2(ALUOut_Out),.SelMux_2(CtrlMux12_2),.Mux_3(CP0_Rdata),.SelMux_3(CtrlMux12_3),.Mux_4(CP1_Rdata),.SelMux_4(CtrlMux12_4),.Mux_5(CountUnit_Out),.SelMux_5(CtrlMux12_5),.Mux_6(Hi_Out),.SelMux_6(CtrlMux12_6),.Mux_7(IMMSEXT_Out),.SelMux_7(CtrlMux12_7),.Mux_8(Lo_Out),.SelMux_8(CtrlMux12_8),.Mux_9(MemDataSel_Out),.SelMux_9(CtrlMux12_9),.Mux_10(PC_Out),.SelMux_10(CtrlMux12_10),.Mux_11({31'b0, LLbit_Out}),.SelMux_11(CtrlMux12_11),.Out(Mux12_Out));
Mux3_5module Mux13(.Mux_1(5'd31),.SelMux_1(CtrlMux13_1),.Mux_2(IR_Out[15:11]),.SelMux_2(CtrlMux13_2),.Mux_3(IR_Out[20:16]),.SelMux_3(CtrlMux13_3),.Out(Mux13_Out));
Mux2_32module Mux14(.Mux_1(GPR_Rdata1),.SelMux_1(CtrlMux14_1),.Mux_2(SEXT_Out),.SelMux_2(CtrlMux14_2),.Out(Mux14_Out));
Mux3_32module Mux15(.Mux_1(GPR_Rdata2),.SelMux_1(CtrlMux15_1),.Mux_2(IMMEXT_Out),.SelMux_2(CtrlMux15_2),.Mux_3(LIMMEXT_Out),.SelMux_3(CtrlMux15_3),.Out(Mux15_Out));
Mux3_32module Mux16(.Mux_1(A_Out),.SelMux_1(CtrlMux16_1),.Mux_2(PC_CIA),.SelMux_2(CtrlMux16_2),.Mux_3(PC_Out),.SelMux_3(CtrlMux16_3),.Out(Mux16_Out));
Mux2_32module Mux17(.Mux_1(B_Out),.SelMux_1(CtrlMux17_1),.Mux_2(SEXT_Out),.SelMux_2(CtrlMux17_2),.Out(Mux17_Out));
Mux9_6module Mux18(.Mux_1(6'b000000),.SelMux_1(CtrlMux18_1),.Mux_2(6'b000001),.SelMux_2(CtrlMux18_2),.Mux_3(6'b000010),.SelMux_3(CtrlMux18_3),.Mux_4(6'b000011),.SelMux_4(CtrlMux18_4),.Mux_5(6'b000110),.SelMux_5(CtrlMux18_5),.Mux_6(6'b000111),.SelMux_6(CtrlMux18_6),.Mux_7(6'b001100),.SelMux_7(CtrlMux18_7),.Mux_8(6'b010010),.SelMux_8(CtrlMux18_8),.Mux_9(6'b010111),.SelMux_9(CtrlMux18_9),.Out(Mux18_Out));
Mux2_32module Mux19(.Mux_1(ALU_Out),.SelMux_1(CtrlMux19_1),.Mux_2(SU_Out),.SelMux_2(CtrlMux19_2),.Out(Mux19_Out));
Mux1_26module Mux20(.Mux_1(IR_Out[25:0]),.SelMux_1(CtrlMux20_1),.Out(Mux20_Out));
Mux1_4module Mux21(.Mux_1(PC_CIA[31:28]),.SelMux_1(CtrlMux21_1),.Out(Mux21_Out));
Mux1_16module Mux22(.Mux_1(IR_Out[15:0]),.SelMux_1(CtrlMux22_1),.Out(Mux22_Out));
Mux1_16module Mux23(.Mux_1(IR_Out[15:0]),.SelMux_1(CtrlMux23_1),.Out(Mux23_Out));
Mux1_16module Mux24(.Mux_1(IR_Out[15:0]),.SelMux_1(CtrlMux24_1),.Out(Mux24_Out));
Mux1_16module Mux25(.Mux_1(IR_Out[15:0]),.SelMux_1(CtrlMux25_1),.Out(Mux25_Out));
Mux2_32module Mux26(.Mux_1(32'b0),.SelMux_1(CtrlMux26_1),.Mux_2(A_Out),.SelMux_2(CtrlMux26_2),.Out(Mux26_Out));
Mux1_32module Mux27(.Mux_1(B_Out),.SelMux_1(CtrlMux27_1),.Out(Mux27_Out));
Mux2_6module Mux28(.Mux_1(6'b000000),.SelMux_1(CtrlMux28_1),.Mux_2(6'b000011),.SelMux_2(CtrlMux28_2),.Out(Mux28_Out));
Mux2_6module Mux29(.Mux_1(6'b000000),.SelMux_1(CtrlMux29_1),.Mux_2(6'b000001),.SelMux_2(CtrlMux29_2),.Out(Mux29_Out));
Mux1_32module Mux30(.Mux_1(A_Out),.SelMux_1(CtrlMux30_1),.Out(Mux30_Out));
Mux3_32module Mux31(.Mux_1(DMem_Out),.SelMux_1(CtrlMux31_1),.Mux_2(GPR_Rdata2),.SelMux_2(CtrlMux31_2),.Mux_3({24'b0,GPR_Rdata2[7:0]}),.SelMux_3(CtrlMux31_3),.Out(Mux31_Out));
Mux1_32module Mux32(.Mux_1(GPR_Rdata2),.SelMux_1(CtrlMux32_1),.Out(Mux32_Out));
Mux2_32module Mux33(.Mux_1(GPR_Rdata1),.SelMux_1(CtrlMux33_1),.Mux_2(MDU_hi),.SelMux_2(CtrlMux33_2),.Out(Mux33_Out));
Mux2_32module Mux34(.Mux_1(GPR_Rdata1),.SelMux_1(CtrlMux34_1),.Mux_2(MDU_lo),.SelMux_2(CtrlMux34_2),.Out(Mux34_Out));
Mux1_1module Mux35(.Mux_1(1'b1),.SelMux_1(CtrlMux35_1),.Out(Mux35_Out));
Mux1_32module Mux36(.Mux_1(A_Out),.SelMux_1(CtrlMux36_1),.Out(Mux36_Out));
Mux1_32module Mux37(.Mux_1(B_Out),.SelMux_1(CtrlMux37_1),.Out(Mux37_Out));
Mux8_6module Mux38(.Mux_1(6'b000001),.SelMux_1(CtrlMux38_1),.Mux_2(6'b000010),.SelMux_2(CtrlMux38_2),.Mux_3(6'b000011),.SelMux_3(CtrlMux38_3),.Mux_4(6'b000100),.SelMux_4(CtrlMux38_4),.Mux_5(6'b000101),.SelMux_5(CtrlMux38_5),.Mux_6(6'b000110),.SelMux_6(CtrlMux38_6),.Mux_7(6'b000111),.SelMux_7(CtrlMux38_7),.Mux_8(6'b001000),.SelMux_8(CtrlMux38_8),.Out(Mux38_Out));
Mux1_32module Mux39(.Mux_1(Hi_Out),.SelMux_1(CtrlMux39_1),.Out(Mux39_Out));
Mux1_32module Mux40(.Mux_1(Lo_Out),.SelMux_1(CtrlMux40_1),.Out(Mux40_Out));
Mux11_6module Mux41(.Mux_1(6'b000001),.SelMux_1(CtrlMux41_1),.Mux_2(6'b000010),.SelMux_2(CtrlMux41_2),.Mux_3(6'b000011),.SelMux_3(CtrlMux41_3),.Mux_4(6'b000100),.SelMux_4(CtrlMux41_4),.Mux_5(6'b000101),.SelMux_5(CtrlMux41_5),.Mux_6(6'b001001),.SelMux_6(CtrlMux41_6),.Mux_7(6'b001010),.SelMux_7(CtrlMux41_7),.Mux_8(6'b010001),.SelMux_8(CtrlMux41_8),.Mux_9(6'b010011),.SelMux_9(CtrlMux41_9),.Mux_10(6'b010100),.SelMux_10(CtrlMux41_10),.Mux_11(6'b010101),.SelMux_11(CtrlMux41_11),.Out(Mux41_Out));
Mux1_2module Mux42(.Mux_1(ALUOut_Out[1:0]),.SelMux_1(CtrlMux42_1),.Out(Mux42_Out));
Mux1_32module Mux43(.Mux_1(DR_Out),.SelMux_1(CtrlMux43_1),.Out(Mux43_Out));
Mux2_32module Mux44(.Mux_1(B_Out),.SelMux_1(CtrlMux44_1),.Mux_2(DR0_Out),.SelMux_2(CtrlMux44_2),.Out(Mux44_Out));
Mux1_1module Mux45(.Mux_1(ALU_OV),.SelMux_1(CtrlMux45_1),.Out(Mux45_Out));
Mux4_1module Mux46(.Mux_1(CMPU_gt),.SelMux_1(CtrlMux46_1),.Mux_2(CMPU_lt),.SelMux_2(CtrlMux46_2),.Mux_3(CMPU_zero),.SelMux_3(CtrlMux46_3),.Mux_4(CP1_fp),.SelMux_4(CtrlMux46_4),.Out(Mux46_Out));
Mux1_8module Mux47(.Mux_1(CP0_ASID),.SelMux_1(CtrlMux47_1),.Out(Mux47_Out));
Mux1_32module Mux48(.Mux_1(B_Out),.SelMux_1(CtrlMux48_1),.Out(Mux48_Out));
Mux3_6module Mux49(.Mux_1(6'b000100),.SelMux_1(CtrlMux49_1),.Mux_2(6'b000101),.SelMux_2(CtrlMux49_2),.Mux_3(6'b000110),.SelMux_3(CtrlMux49_3),.Out(Mux49_Out));
Mux2_5module Mux50(.Mux_1(A_Out[4:0]),.SelMux_1(CtrlMux50_1),.Mux_2(IR_Out[10:6]),.SelMux_2(CtrlMux50_2),.Out(Mux50_Out));
Mux2_8module Mux51(.Mux_1(8'd0),.SelMux_1(CtrlMux51_1),.Mux_2(PIDReg_Out),.SelMux_2(CtrlMux51_2),.Out(Mux51_Out));
Mux1_32module Mux52(.Mux_1(PC_Out),.SelMux_1(CtrlMux52_1),.Out(Mux52_Out));
Mux2_5module Mux53(.Mux_1(5'h08),.SelMux_1(CtrlMux53_1),.Mux_2(5'h0d),.SelMux_2(CtrlMux53_2),.Out(Mux53_Out));
Mux1_5module Mux54(.Mux_1(IR_Out[15:11]),.SelMux_1(CtrlMux54_1),.Out(Mux54_Out));
Mux1_32module Mux55(.Mux_1(A_Out),.SelMux_1(CtrlMux55_1),.Out(Mux55_Out));
Mux1_5module Mux56(.Mux_1(IR_Out[15:11]),.SelMux_1(CtrlMux56_1),.Out(Mux56_Out));
Mux1_3module Mux57(.Mux_1(IR_Out[20:18]),.SelMux_1(CtrlMux57_1),.Out(Mux57_Out));
Mux1_5module Mux58(.Mux_1(IR_Out[15:11]),.SelMux_1(CtrlMux58_1),.Out(Mux58_Out));
Mux1_1module Mux59(.Mux_1(IR_Out[16]),.SelMux_1(CtrlMux59_1),.Out(Mux59_Out));
Mux1_32module Mux60(.Mux_1(A_Out),.SelMux_1(CtrlMux60_1),.Out(Mux60_Out));
Mux1_5module Mux61(.Mux_1(IR_Out[15:11]),.SelMux_1(CtrlMux61_1),.Out(Mux61_Out));
Mux1_1module Mux64(.Mux_1(ConditionReg_Out),.SelMux_1(CtrlMux64_1),.Out(Mux64_Out));
Mux1_1module Mux65(.Mux_1(ConditionReg_Out),.SelMux_1(CtrlMux65_1),.Out(Mux65_Out));
Mux1_32module Mux68(.Mux_1(IR_Out),.SelMux_1(CtrlMux68_1),.Out(Mux68_Out));
Mux1_1module Mux69(.Mux_1(LLbit_Out),.SelMux_1(CtrlMux69_1),.Out(Mux69_Out));
Mux1_1module Mux70(.Mux_1(ConditionReg_Out),.SelMux_1(CtrlMux70_1),.Out(Mux70_Out));
Mux1_1module Mux71(.Mux_1(OVReg_Out),.SelMux_1(CtrlMux71_1),.Out(Mux71_Out));
Mux1_1module Mux72(.Mux_1(ConditionReg_Out),.SelMux_1(CtrlMux72_1),.Out(Mux72_Out));
endmodule
