module CPU(clr,clk);
input clk,clr;
wire CtrlMux2_1;
wire [31:0]Mux2_Out;
wire CtrlMux3_1;
wire [31:0]Mux3_Out;
wire CtrlMux8_1;
wire [31:0]Mux8_Out;
wire CtrlMux9_1;
wire [4:0]Mux9_Out;
wire CtrlMux10_1;
wire [4:0]Mux10_Out;
wire CtrlMux11_1;
wire [31:0]Mux11_Out;
wire CtrlMux12_1;
wire [4:0]Mux12_Out;
wire CtrlMux13_1;
wire [31:0]Mux13_Out;
wire CtrlMux14_1;
wire [31:0]Mux14_Out;
wire CtrlMux15_1;
wire [31:0]Mux15_Out;
wire CtrlMux16_1;
wire [31:0]Mux16_Out;
wire CtrlMux17_1;
wire [5:0]Mux17_Out;
wire CtrlMux18_1;
wire [31:0]Mux18_Out;
wire CtrlMux42_1;
wire Mux42_Out;
wire CtrlMux65_1;
wire [5:0]Mux65_Out;
wire CtrlMux68_1;
wire Mux68_Out;
wire [5:0]CU_Func;
wire CtrlPCInc;
wire [31:0]PC_Out;
wire [31:0]IMem_Out;
wire CtrlIR;
wire [31:0]IR_Out;
wire CtrlRegs;
wire [31:0]Regs_Rdata1;
wire [31:0]Regs_Rdata2;
wire CtrlA;
wire [31:0]A_Out;
wire CtrlB;
wire [31:0]B_Out;
wire CtrlALUOut;
wire [31:0]ALUOut_Out;
wire [31:0]ALU_Out;
wire ALU_OV;
wire [31:0]CP0_ASID;
wire CtrlOVReg;
wire OVReg_Out;
CU_module CU(.clr(clr),.clk(clk),.Op(IR_Out[31:26]),.IRFunc(Mux65_Out),.OV(Mux68_Out),.Func(CU_Func),.CtrlA(CtrlA),.CtrlALUOut(CtrlALUOut),.CtrlB(CtrlB),.CtrlIR(CtrlIR),.CtrlOVReg(CtrlOVReg),.CtrlPCInc(CtrlPCInc),.CtrlRegs(CtrlRegs),.CtrlMux2_1(CtrlMux2_1),.CtrlMux3_1(CtrlMux3_1),.CtrlMux8_1(CtrlMux8_1),.CtrlMux9_1(CtrlMux9_1),.CtrlMux10_1(CtrlMux10_1),.CtrlMux11_1(CtrlMux11_1),.CtrlMux12_1(CtrlMux12_1),.CtrlMux13_1(CtrlMux13_1),.CtrlMux14_1(CtrlMux14_1),.CtrlMux15_1(CtrlMux15_1),.CtrlMux16_1(CtrlMux16_1),.CtrlMux17_1(CtrlMux17_1),.CtrlMux18_1(CtrlMux18_1),.CtrlMux42_1(CtrlMux42_1),.CtrlMux65_1(CtrlMux65_1),.CtrlMux68_1(CtrlMux68_1));
PC_module PC(.clr(clr),.CtrlPCInc(CtrlPCInc),.Out(PC_Out));
IMemory_module IMem(.clr(clr),.RAddr(Mux3_Out),.ASID(Mux2_Out),.Out(IMem_Out));
IR_module IR(.clr(clr),.In(Mux8_Out),.CtrlIR(CtrlIR),.Out(IR_Out));
Regs_module Regs(.clr(clr),.CtrlRegs(CtrlRegs),.RReg1(Mux9_Out),.RReg2(Mux10_Out),.WReg(Mux12_Out),.WData(Mux11_Out),.Rdata1(Regs_Rdata1),.Rdata2(Regs_Rdata2));
A_module A(.clr(clr),.CtrlA(CtrlA),.In(Mux13_Out),.Out(A_Out));
B_module B(.clr(clr),.CtrlB(CtrlB),.In(Mux14_Out),.Out(B_Out));
ALUOut_module ALUOut(.clr(clr),.CtrlALUOut(CtrlALUOut),.In(Mux18_Out),.Out(ALUOut_Out));
ALU_module ALU(.A(Mux15_Out),.B(Mux16_Out),.Func(Mux17_Out),.Out(ALU_Out),.OV(ALU_OV));
CP0_module CP0(.clr(clr),.ASID(CP0_ASID));
OVReg_module OVReg(.clr(clr),.CtrlOVReg(CtrlOVReg),.In(Mux42_Out),.Out(OVReg_Out));
Mux1_32module Mux2(.Mux_1(CP0_ASID),.SelMux_1(CtrlMux2_1),.Out(Mux2_Out));
Mux1_32module Mux3(.Mux_1(PC_Out),.SelMux_1(CtrlMux3_1),.Out(Mux3_Out));
Mux1_32module Mux8(.Mux_1(IMem_Out),.SelMux_1(CtrlMux8_1),.Out(Mux8_Out));
Mux1_5module Mux9(.Mux_1(IR_Out[25:21]),.SelMux_1(CtrlMux9_1),.Out(Mux9_Out));
Mux1_5module Mux10(.Mux_1(IR_Out[20:16]),.SelMux_1(CtrlMux10_1),.Out(Mux10_Out));
Mux1_32module Mux11(.Mux_1(ALUOut_Out),.SelMux_1(CtrlMux11_1),.Out(Mux11_Out));
Mux1_5module Mux12(.Mux_1(IR_Out[15:11]),.SelMux_1(CtrlMux12_1),.Out(Mux12_Out));
Mux1_32module Mux13(.Mux_1(Regs_Rdata1),.SelMux_1(CtrlMux13_1),.Out(Mux13_Out));
Mux1_32module Mux14(.Mux_1(Regs_Rdata2),.SelMux_1(CtrlMux14_1),.Out(Mux14_Out));
Mux1_32module Mux15(.Mux_1(A_Out),.SelMux_1(CtrlMux15_1),.Out(Mux15_Out));
Mux1_32module Mux16(.Mux_1(B_Out),.SelMux_1(CtrlMux16_1),.Out(Mux16_Out));
Mux1_6module Mux17(.Mux_1(CU_Func),.SelMux_1(CtrlMux17_1),.Out(Mux17_Out));
Mux1_32module Mux18(.Mux_1(ALU_Out),.SelMux_1(CtrlMux18_1),.Out(Mux18_Out));
Mux1_1module Mux42(.Mux_1(ALU_OV),.SelMux_1(CtrlMux42_1),.Out(Mux42_Out));
Mux1_6module Mux65(.Mux_1(IR_Out[5:0]),.SelMux_1(CtrlMux65_1),.Out(Mux65_Out));
Mux1_1module Mux68(.Mux_1(OVReg_Out),.SelMux_1(CtrlMux68_1),.Out(Mux68_Out));
endmodule
