module CU_module(clr,clk,Op,IRFunc,OV,Func,CtrlA,CtrlALUOut,CtrlB,CtrlIR,CtrlOVReg,CtrlPCInc,CtrlRegs,CtrlMux2_1,CtrlMux3_1,CtrlMux8_1,CtrlMux9_1,CtrlMux10_1,CtrlMux11_1,CtrlMux12_1,CtrlMux13_1,CtrlMux14_1,CtrlMux15_1,CtrlMux16_1,CtrlMux17_1,CtrlMux18_1,CtrlMux42_1,CtrlMux65_1,CtrlMux68_1);
input clr;
input clk;
input [5:0]Op;
input [5:0]IRFunc;
input OV;
output [5:0]Func;
output CtrlA;
output CtrlALUOut;
output CtrlB;
output CtrlIR;
output CtrlOVReg;
output CtrlPCInc;
output CtrlRegs;
output CtrlMux2_1;
output CtrlMux3_1;
output CtrlMux8_1;
output CtrlMux9_1;
output CtrlMux10_1;
output CtrlMux11_1;
output CtrlMux12_1;
output CtrlMux13_1;
output CtrlMux14_1;
output CtrlMux15_1;
output CtrlMux16_1;
output CtrlMux17_1;
output CtrlMux18_1;
output CtrlMux42_1;
output CtrlMux65_1;
output CtrlMux68_1;
wire P0,P1,P2,P3,P4,P;
wire IRFunc22;
wire OP00;
Initial_model Initial(.clr(clr),.clk(clk),.P0(P0),.P1(P1),.P2(P2),.P3(P3),.P4(P4),.P(P),.Op(Op),.IRFunc(IRFunc),.Func(Func),.IRFunc22(IRFunc22),.OP00(OP00));
assign CtrlA=(P1&OP00&IRFunc22);
assign CtrlALUOut=(P2&OP00&IRFunc22);
assign CtrlB=(P1&OP00&IRFunc22);
assign CtrlIR=(P0&OP00&IRFunc22);
assign CtrlMux10_1=(P0&OP00&IRFunc22);
assign CtrlMux11_1=(P3&OP00&IRFunc22);
assign CtrlMux12_1=(P3&OP00&IRFunc22);
assign CtrlMux13_1=(P0&OP00&IRFunc22);
assign CtrlMux14_1=(P0&OP00&IRFunc22);
assign CtrlMux15_1=(P1&OP00&IRFunc22);
assign CtrlMux16_1=(P1&OP00&IRFunc22);
assign CtrlMux17_1=(P1&OP00&IRFunc22);
assign CtrlMux18_1=(P1&OP00&IRFunc22);
assign CtrlMux2_1=((P|P5));
assign CtrlMux3_1=((P|P5));
assign CtrlMux42_1=(P1&OP00&IRFunc22);
assign CtrlMux65_1=(P0&OP00&IRFunc22);
assign CtrlMux68_1=(P3&OP00&IRFunc22);
assign CtrlMux8_1=((P|P5));
assign CtrlMux9_1=(P0&OP00&IRFunc22);
assign CtrlOVReg=(P2&OP00&IRFunc22);
assign CtrlPCInc=(P0&OP00&IRFunc22);
assign CtrlRegs=(P4&OP00&IRFunc22);
endmodule
